/* Automatically generated from https://wokwi.com/projects/376553022662786049 */

`default_nettype none

module tt_um_wokwi_376553022662786049(
  input  wire [7:0] ui_in,    // Dedicated inputs
  output wire [7:0] uo_out,    // Dedicated outputs
  input  wire [7:0] uio_in,    // IOs: Input path
  output wire [7:0] uio_out,    // IOs: Output path
  output wire [7:0] uio_oe,    // IOs: Enable path (active high: 0=input, 1=output)
  input ena,
  input clk,
  input rst_n
);
  wire net1 = clk;
  wire net2 = ui_in[0];
  wire net3 = ui_in[1];
  wire net4 = ui_in[2];
  wire net5 = ui_in[3];
  wire net6 = ui_in[4];
  wire net7 = ui_in[5];
  wire net8 = ui_in[6];
  wire net9 = ui_in[7];
  wire net10;
  wire net11;
  wire net12;
  wire net13;
  wire net14;
  wire net15;
  wire net16;
  wire net17;
  wire net18 = 1'b1;
  wire net19;
  wire net20 = 1'b1;
  wire net21;
  wire net22 = 1'b1;
  wire net23;
  wire net24 = 1'b1;
  wire net25;
  wire net26 = 1'b1;
  wire net27 = uio_in[5];
  wire net28 = 1'b0;
  wire net29 = uio_in[6];
  wire net30 = 1'b0;
  wire net31;
  wire net32 = 1'b1;
  wire net33 = 1'b1;
  wire net34 = 1'b0;
  wire net35 = 1'b0;
  wire net36 = 1'b0;
  wire net37;
  wire net38;
  wire net39;
  wire net40;
  wire net41;
  wire net42 = 1'b0;
  wire net43;
  wire net44;
  wire net45;
  wire net46;
  wire net47;
  wire net48;
  wire net49;
  wire net50;
  wire net51;
  wire net52;
  wire net53;
  wire net54;
  wire net55;
  wire net56;
  wire net57;
  wire net58;
  wire net59 = 1'b0;
  wire net60;
  wire net61;
  wire net62;
  wire net63;
  wire net64;
  wire net65;
  wire net66;
  wire net67;
  wire net68;
  wire net69;
  wire net70;
  wire net71;
  wire net72 = 1'b0;
  wire net73;
  wire net74 = 1'b0;
  wire net75;
  wire net76;
  wire net77;
  wire net78;
  wire net79;
  wire net80;
  wire net81;
  wire net82;
  wire net83;
  wire net84 = 1'b0;
  wire net85;
  wire net86 = 1'b0;
  wire net87;
  wire net88;
  wire net89;
  wire net90;
  wire net91;
  wire net92;
  wire net93 = 1'b0;
  wire net94;
  wire net95 = 1'b0;
  wire net96;
  wire net97;
  wire net98;
  wire net99 = 1'b0;
  wire net100;
  wire net101 = 1'b0;
  wire net102;
  wire net103;
  wire net104;
  wire net105;
  wire net106;
  wire net107;
  wire net108;
  wire net109;
  wire net110;
  wire net111;
  wire net112;
  wire net113;
  wire net114;
  wire net115 = 1'b0;
  wire net116;
  wire net117 = 1'b0;
  wire net118;
  wire net119;
  wire net120;
  wire net121;
  wire net122;
  wire net123;
  wire net124;
  wire net125;
  wire net126;
  wire net127;
  wire net128;
  wire net129;
  wire net130;
  wire net131 = 1'b0;
  wire net132;
  wire net133 = 1'b0;
  wire net134;
  wire net135;
  wire net136;
  wire net137;
  wire net138;
  wire net139;
  wire net140;
  wire net141;
  wire net142;
  wire net143;
  wire net144;
  wire net145;
  wire net146;
  wire net147 = 1'b0;
  wire net148;
  wire net149 = 1'b0;
  wire net150;
  wire net151;
  wire net152;
  wire net153;
  wire net154;
  wire net155;
  wire net156;
  wire net157;
  wire net158;
  wire net159;
  wire net160;
  wire net161;
  wire net162;
  wire net163 = 1'b0;
  wire net164;
  wire net165 = 1'b0;
  wire net166;
  wire net167;
  wire net168;
  wire net169;
  wire net170;
  wire net171;
  wire net172;
  wire net173;
  wire net174;
  wire net175;
  wire net176;
  wire net177;
  wire net178;
  wire net179 = 1'b0;
  wire net180;
  wire net181 = 1'b0;
  wire net182;
  wire net183;
  wire net184;
  wire net185;
  wire net186;
  wire net187;
  wire net188;
  wire net189;
  wire net190;
  wire net191;
  wire net192;
  wire net193;
  wire net194;
  wire net195 = 1'b0;
  wire net196;
  wire net197 = 1'b0;
  wire net198;
  wire net199;
  wire net200;
  wire net201;
  wire net202;
  wire net203;
  wire net204;
  wire net205;
  wire net206;
  wire net207;
  wire net208;
  wire net209;
  wire net210;
  wire net211 = 1'b0;
  wire net212;
  wire net213 = 1'b0;
  wire net214;
  wire net215;
  wire net216;
  wire net217;
  wire net218;
  wire net219;
  wire net220;
  wire net221;
  wire net222;
  wire net223;
  wire net224;
  wire net225;
  wire net226;
  wire net227 = 1'b0;
  wire net228;
  wire net229 = 1'b0;
  wire net230;
  wire net231;
  wire net232;
  wire net233;
  wire net234;
  wire net235;
  wire net236;
  wire net237;
  wire net238;
  wire net239;
  wire net240;
  wire net241;
  wire net242;
  wire net243 = 1'b0;
  wire net244;
  wire net245 = 1'b0;
  wire net246;
  wire net247;
  wire net248;
  wire net249;
  wire net250;
  wire net251;
  wire net252;
  wire net253;
  wire net254;
  wire net255;
  wire net256;
  wire net257;
  wire net258;
  wire net259 = 1'b0;
  wire net260 = 1'b0;
  wire net261;
  wire net262;
  wire net263;
  wire net264;
  wire net265 = 1'b0;
  wire net266;
  wire net267;
  wire net268;
  wire net269;
  wire net270 = 1'b0;
  wire net271;
  wire net272 = 1'b0;
  wire net273;
  wire net274;
  wire net275;
  wire net276;
  wire net277 = 1'b0;
  wire net278;
  wire net279 = 1'b0;
  wire net280;
  wire net281;
  wire net282;
  wire net283;
  wire net284 = 1'b0;
  wire net285;
  wire net286 = 1'b0;
  wire net287;
  wire net288;
  wire net289;
  wire net290;
  wire net291 = 1'b0;
  wire net292;
  wire net293 = 1'b0;
  wire net294;
  wire net295;
  wire net296;
  wire net297;
  wire net298 = 1'b0;
  wire net299;
  wire net300 = 1'b0;
  wire net301;
  wire net302;
  wire net303;
  wire net304;
  wire net305;
  wire net306;
  wire net307;
  wire net308 = 1'b0;
  wire net309;
  wire net310 = 1'b0;
  wire net311;
  wire net312;
  wire net313;
  wire net314;
  wire net315 = 1'b0;
  wire net316;
  wire net317;
  wire net318 = 1'b0;
  wire net319;
  wire net320;
  wire net321;
  wire net322;
  wire net323 = 1'b0;
  wire net324;
  wire net325 = 1'b0;
  wire net326;
  wire net327;
  wire net328;
  wire net329;
  wire net330;
  wire net331;
  wire net332;
  wire net333 = 1'b0;
  wire net334 = 1'b0;
  wire net335;
  wire net336 = 1'b0;
  wire net337;
  wire net338;
  wire net339;
  wire net340;
  wire net341 = 1'b0;
  wire net342;
  wire net343 = 1'b0;
  wire net344;
  wire net345;
  wire net346;
  wire net347;
  wire net348;
  wire net349;
  wire net350;
  wire net351 = 1'b0;
  wire net352;
  wire net353 = 1'b0;
  wire net354;
  wire net355;
  wire net356;
  wire net357;
  wire net358 = 1'b0;
  wire net359;
  wire net360 = 1'b0;
  wire net361;
  wire net362;
  wire net363;
  wire net364;
  wire net365;
  wire net366;
  wire net367;
  wire net368 = 1'b0;
  wire net369;
  wire net370 = 1'b0;
  wire net371;
  wire net372;
  wire net373;
  wire net374;
  wire net375 = 1'b0;
  wire net376;
  wire net377 = 1'b0;
  wire net378;
  wire net379;
  wire net380;
  wire net381;
  wire net382;
  wire net383;
  wire net384;
  wire net385 = 1'b0;
  wire net386;
  wire net387;
  wire net388 = 1'b0;
  wire net389;
  wire net390;
  wire net391;
  wire net392;
  wire net393;
  wire net394;
  wire net395;
  wire net396;
  wire net397;
  wire net398;
  wire net399;
  wire net400;
  wire net401;
  wire net402;
  wire net403;
  wire net404;
  wire net405;
  wire net406;
  wire net407 = 1'b0;
  wire net408;
  wire net409;
  wire net410;
  wire net411;
  wire net412;
  wire net413;
  wire net414;
  wire net415;
  wire net416;
  wire net417;
  wire net418;
  wire net419;
  wire net420;
  wire net421 = 1'b0;
  wire net422;
  wire net423 = 1'b0;
  wire net424;
  wire net425;
  wire net426;
  wire net427;
  wire net428;
  wire net429;
  wire net430;
  wire net431 = 1'b0;
  wire net432;
  wire net433 = 1'b0;
  wire net434;
  wire net435;
  wire net436;
  wire net437;
  wire net438;
  wire net439;
  wire net440;
  wire net441;
  wire net442;
  wire net443;
  wire net444;
  wire net445;
  wire net446;
  wire net447 = 1'b0;
  wire net448;
  wire net449 = 1'b0;
  wire net450;
  wire net451;
  wire net452;
  wire net453;
  wire net454;
  wire net455;
  wire net456;
  wire net457 = 1'b0;
  wire net458;
  wire net459 = 1'b0;
  wire net460;
  wire net461;
  wire net462;
  wire net463;
  wire net464;
  wire net465;
  wire net466;
  wire net467;
  wire net468;
  wire net469;
  wire net470;
  wire net471;
  wire net472;
  wire net473 = 1'b0;
  wire net474;
  wire net475 = 1'b0;
  wire net476;
  wire net477;
  wire net478;
  wire net479;
  wire net480;
  wire net481;
  wire net482;
  wire net483 = 1'b0;
  wire net484;
  wire net485 = 1'b0;
  wire net486;
  wire net487;
  wire net488;
  wire net489;
  wire net490;
  wire net491;
  wire net492;
  wire net493;
  wire net494;
  wire net495;
  wire net496;
  wire net497;
  wire net498;
  wire net499 = 1'b0;
  wire net500;
  wire net501 = 1'b0;
  wire net502;
  wire net503;
  wire net504;
  wire net505 = 1'b0;
  wire net506;
  wire net507 = 1'b0;
  wire net508;
  wire net509;
  wire net510;
  wire net511;
  wire net512;
  wire net513;
  wire net514 = 1'b0;
  wire net515 = 1'b0;
  wire net516;
  wire net517;
  wire net518 = 1'b0;
  wire net519;
  wire net520;
  wire net521;
  wire net522;
  wire net523;
  wire net524;
  wire net525;
  wire net526 = 1'b0;
  wire net527;
  wire net528;
  wire net529 = 1'b0;
  wire net530;
  wire net531;
  wire net532;
  wire net533;
  wire net534;
  wire net535;
  wire net536;
  wire net537 = 1'b0;
  wire net538 = 1'b0;
  wire net539;
  wire net540;
  wire net541;
  wire net542;
  wire net543;
  wire net544;
  wire net545;
  wire net546 = 1'b0;
  wire net547;
  wire net548 = 1'b0;
  wire net549;
  wire net550;
  wire net551;
  wire net552;
  wire net553;
  wire net554;
  wire net555;
  wire net556 = 1'b0;
  wire net557;
  wire net558 = 1'b0;
  wire net559;
  wire net560;
  wire net561;
  wire net562;
  wire net563;
  wire net564;
  wire net565;
  wire net566 = 1'b0;
  wire net567;
  wire net568;
  wire net569 = 1'b0;
  wire net570;
  wire net571;
  wire net572;
  wire net573;
  wire net574;
  wire net575;
  wire net576;
  wire net577 = 1'b0;
  wire net578;
  wire net579;
  wire net580 = 1'b0;
  wire net581;
  wire net582;
  wire net583;
  wire net584;
  wire net585;
  wire net586;
  wire net587;
  wire net588 = 1'b0;

  assign uo_out[0] = net1;
  assign uo_out[1] = net10;
  assign uo_out[2] = net11;
  assign uo_out[3] = net12;
  assign uo_out[4] = net13;
  assign uo_out[5] = net14;
  assign uo_out[6] = net15;
  assign uo_out[7] = net16;
  assign uio_out[0] = net17;
  assign uio_oe[0] = net18;
  assign uio_out[1] = net19;
  assign uio_oe[1] = net20;
  assign uio_out[2] = net21;
  assign uio_oe[2] = net22;
  assign uio_out[3] = net23;
  assign uio_oe[3] = net24;
  assign uio_out[4] = net25;
  assign uio_oe[4] = net26;
  assign uio_out[5] = net28;
  assign uio_oe[5] = net28;
  assign uio_out[6] = net30;
  assign uio_oe[6] = net30;
  assign uio_out[7] = net31;
  assign uio_oe[7] = net32;

  dff_cell flop1 (
    .d (net37),
    .clk (net1),
    .q (net38)
  );
  dff_cell flop2 (
    .d (net38),
    .clk (net1),
    .q (net39)
  );
  dff_cell flop3 (
    .d (net39),
    .clk (net1),
    .q (net40)
  );
  dff_cell flop4 (
    .d (net40),
    .clk (net1),
    .q (net10)
  );
  xor_cell xor3 (
    .a (net10),
    .b (net40),
    .out (net37)
  );
  dffsr_cell flop28 (
    .d (net41),
    .clk (net16),
    .s (net42),
    .r (net42),
    .q (net43),
    .notq (net41)
  );
  dffsr_cell flop29 (
    .d (net44),
    .clk (net41),
    .s (net42),
    .r (net42),
    .q (net45),
    .notq (net44)
  );
  dffsr_cell flop30 (
    .d (net46),
    .clk (net44),
    .s (net42),
    .r (net42),
    .q (net47),
    .notq (net46)
  );
  dffsr_cell flop31 (
    .d (net48),
    .clk (net46),
    .s (net42),
    .r (net42),
    .q (net49),
    .notq (net48)
  );
  dffsr_cell flop32 (
    .d (net50),
    .clk (net48),
    .s (net42),
    .r (net42),
    .q (net51),
    .notq (net50)
  );
  dffsr_cell flop33 (
    .d (net52),
    .clk (net50),
    .s (net42),
    .r (net42),
    .q (net53),
    .notq (net52)
  );
  and_cell and21 (
    .a (net43),
    .b (net45),
    .out (net54)
  );
  and_cell and22 (
    .a (net54),
    .b (net47),
    .out (net55)
  );
  and_cell and23 (
    .a (net55),
    .b (net56),
    .out (net15)
  );
  and_cell and24 (
    .a (net49),
    .b (net51),
    .out (net57)
  );
  and_cell and25 (
    .a (net57),
    .b (net53),
    .out (net56)
  );
  dffsr_cell flop20 (
    .d (net58),
    .clk (net16),
    .s (net59),
    .r (net59),
    .q (net60),
    .notq (net58)
  );
  dffsr_cell flop21 (
    .d (net61),
    .clk (net58),
    .s (net59),
    .r (net59),
    .q (net62),
    .notq (net61)
  );
  dffsr_cell flop22 (
    .d (net63),
    .clk (net61),
    .s (net59),
    .r (net59),
    .q (net64),
    .notq (net63)
  );
  dffsr_cell flop24 (
    .d (net65),
    .clk (net63),
    .s (net59),
    .r (net59),
    .q (net66),
    .notq (net65)
  );
  dffsr_cell flop25 (
    .d (net67),
    .clk (net65),
    .s (net59),
    .r (net59),
    .q (net68),
    .notq (net67)
  );
  and_cell and10 (
    .a (net60),
    .b (net62),
    .out (net69)
  );
  and_cell and11 (
    .a (net69),
    .b (net64),
    .out (net70)
  );
  and_cell and12 (
    .a (net70),
    .b (net66),
    .out (net71)
  );
  and_cell and13 (
    .a (net71),
    .b (net68),
    .out (net14)
  );
  dffsr_cell flop26 (
    .d (net73),
    .clk (net16),
    .s (net74),
    .r (net74),
    .q (net75),
    .notq (net73)
  );
  dffsr_cell flop27 (
    .d (net76),
    .clk (net73),
    .s (net74),
    .r (net74),
    .q (net77),
    .notq (net76)
  );
  dffsr_cell flop34 (
    .d (net78),
    .clk (net76),
    .s (net74),
    .r (net74),
    .q (net79),
    .notq (net78)
  );
  dffsr_cell flop35 (
    .d (net80),
    .clk (net78),
    .s (net74),
    .r (net74),
    .q (net81),
    .notq (net80)
  );
  and_cell and14 (
    .a (net75),
    .b (net77),
    .out (net82)
  );
  and_cell and15 (
    .a (net82),
    .b (net79),
    .out (net83)
  );
  and_cell and16 (
    .a (net83),
    .b (net81),
    .out (net13)
  );
  dffsr_cell flop16 (
    .d (net85),
    .clk (net16),
    .s (net86),
    .r (net86),
    .q (net87),
    .notq (net85)
  );
  dffsr_cell flop17 (
    .d (net88),
    .clk (net85),
    .s (net86),
    .r (net86),
    .q (net89),
    .notq (net88)
  );
  dffsr_cell flop18 (
    .d (net90),
    .clk (net88),
    .s (net86),
    .r (net86),
    .q (net91),
    .notq (net90)
  );
  and_cell and2 (
    .a (net87),
    .b (net89),
    .out (net92)
  );
  and_cell and4 (
    .a (net92),
    .b (net91),
    .out (net12)
  );
  dffsr_cell flop19 (
    .d (net94),
    .clk (net16),
    .s (net95),
    .r (net95),
    .q (net96),
    .notq (net94)
  );
  dffsr_cell flop23 (
    .d (net97),
    .clk (net94),
    .s (net95),
    .r (net95),
    .q (net98),
    .notq (net97)
  );
  and_cell and17 (
    .a (net96),
    .b (net98),
    .out (net11)
  );
  dff_cell flop40 (
    .d (net2),
    .clk (net1),
    .q (net17)
  );
  dffsr_cell flop41 (
    .d (net100),
    .clk (net1),
    .s (net101),
    .r (net101),
    .q (net102),
    .notq (net100)
  );
  dffsr_cell flop42 (
    .d (net103),
    .clk (net100),
    .s (net101),
    .r (net101),
    .q (net104),
    .notq (net103)
  );
  dffsr_cell flop43 (
    .d (net105),
    .clk (net103),
    .s (net101),
    .r (net101),
    .q (net106),
    .notq (net105)
  );
  dffsr_cell flop44 (
    .d (net107),
    .clk (net105),
    .s (net101),
    .r (net101),
    .q (net108),
    .notq (net107)
  );
  dffsr_cell flop45 (
    .d (net109),
    .clk (net107),
    .s (net101),
    .r (net101),
    .q (net110),
    .notq (net109)
  );
  and_cell and18 (
    .a (net102),
    .b (net104),
    .out (net111)
  );
  and_cell and19 (
    .a (net111),
    .b (net106),
    .out (net112)
  );
  and_cell and20 (
    .a (net112),
    .b (net108),
    .out (net113)
  );
  and_cell and35 (
    .a (net113),
    .b (net110),
    .out (net114)
  );
  dffsr_cell flop46 (
    .d (net116),
    .clk (net1),
    .s (net117),
    .r (net117),
    .q (net118),
    .notq (net116)
  );
  dffsr_cell flop47 (
    .d (net119),
    .clk (net116),
    .s (net117),
    .r (net117),
    .q (net120),
    .notq (net119)
  );
  dffsr_cell flop48 (
    .d (net121),
    .clk (net119),
    .s (net117),
    .r (net117),
    .q (net122),
    .notq (net121)
  );
  dffsr_cell flop49 (
    .d (net123),
    .clk (net121),
    .s (net117),
    .r (net117),
    .q (net124),
    .notq (net123)
  );
  dffsr_cell flop50 (
    .d (net125),
    .clk (net123),
    .s (net117),
    .r (net117),
    .q (net126),
    .notq (net125)
  );
  and_cell and36 (
    .a (net118),
    .b (net120),
    .out (net127)
  );
  and_cell and37 (
    .a (net127),
    .b (net122),
    .out (net128)
  );
  and_cell and38 (
    .a (net128),
    .b (net124),
    .out (net129)
  );
  and_cell and39 (
    .a (net129),
    .b (net126),
    .out (net130)
  );
  dffsr_cell flop51 (
    .d (net132),
    .clk (net1),
    .s (net133),
    .r (net133),
    .q (net134),
    .notq (net132)
  );
  dffsr_cell flop52 (
    .d (net135),
    .clk (net132),
    .s (net133),
    .r (net133),
    .q (net136),
    .notq (net135)
  );
  dffsr_cell flop53 (
    .d (net137),
    .clk (net135),
    .s (net133),
    .r (net133),
    .q (net138),
    .notq (net137)
  );
  dffsr_cell flop54 (
    .d (net139),
    .clk (net137),
    .s (net133),
    .r (net133),
    .q (net140),
    .notq (net139)
  );
  dffsr_cell flop55 (
    .d (net141),
    .clk (net139),
    .s (net133),
    .r (net133),
    .q (net142),
    .notq (net141)
  );
  and_cell and40 (
    .a (net134),
    .b (net136),
    .out (net143)
  );
  and_cell and41 (
    .a (net143),
    .b (net138),
    .out (net144)
  );
  and_cell and42 (
    .a (net144),
    .b (net140),
    .out (net145)
  );
  and_cell and43 (
    .a (net145),
    .b (net142),
    .out (net146)
  );
  dffsr_cell flop56 (
    .d (net148),
    .clk (net1),
    .s (net149),
    .r (net149),
    .q (net150),
    .notq (net148)
  );
  dffsr_cell flop57 (
    .d (net151),
    .clk (net148),
    .s (net149),
    .r (net149),
    .q (net152),
    .notq (net151)
  );
  dffsr_cell flop58 (
    .d (net153),
    .clk (net151),
    .s (net149),
    .r (net149),
    .q (net154),
    .notq (net153)
  );
  dffsr_cell flop59 (
    .d (net155),
    .clk (net153),
    .s (net149),
    .r (net149),
    .q (net156),
    .notq (net155)
  );
  dffsr_cell flop60 (
    .d (net157),
    .clk (net155),
    .s (net149),
    .r (net149),
    .q (net158),
    .notq (net157)
  );
  and_cell and44 (
    .a (net150),
    .b (net152),
    .out (net159)
  );
  and_cell and45 (
    .a (net159),
    .b (net154),
    .out (net160)
  );
  and_cell and46 (
    .a (net160),
    .b (net156),
    .out (net161)
  );
  and_cell and47 (
    .a (net161),
    .b (net158),
    .out (net162)
  );
  dffsr_cell flop61 (
    .d (net164),
    .clk (net114),
    .s (net165),
    .r (net165),
    .q (net166),
    .notq (net164)
  );
  dffsr_cell flop62 (
    .d (net167),
    .clk (net164),
    .s (net165),
    .r (net165),
    .q (net168),
    .notq (net167)
  );
  dffsr_cell flop63 (
    .d (net169),
    .clk (net167),
    .s (net165),
    .r (net165),
    .q (net170),
    .notq (net169)
  );
  dffsr_cell flop64 (
    .d (net171),
    .clk (net169),
    .s (net165),
    .r (net165),
    .q (net172),
    .notq (net171)
  );
  dffsr_cell flop65 (
    .d (net173),
    .clk (net171),
    .s (net165),
    .r (net165),
    .q (net174),
    .notq (net173)
  );
  and_cell and48 (
    .a (net166),
    .b (net168),
    .out (net175)
  );
  and_cell and49 (
    .a (net175),
    .b (net170),
    .out (net176)
  );
  and_cell and50 (
    .a (net176),
    .b (net172),
    .out (net177)
  );
  and_cell and51 (
    .a (net177),
    .b (net174),
    .out (net178)
  );
  dffsr_cell flop66 (
    .d (net180),
    .clk (net130),
    .s (net181),
    .r (net181),
    .q (net182),
    .notq (net180)
  );
  dffsr_cell flop67 (
    .d (net183),
    .clk (net180),
    .s (net181),
    .r (net181),
    .q (net184),
    .notq (net183)
  );
  dffsr_cell flop68 (
    .d (net185),
    .clk (net183),
    .s (net181),
    .r (net181),
    .q (net186),
    .notq (net185)
  );
  dffsr_cell flop69 (
    .d (net187),
    .clk (net185),
    .s (net181),
    .r (net181),
    .q (net188),
    .notq (net187)
  );
  dffsr_cell flop70 (
    .d (net189),
    .clk (net187),
    .s (net181),
    .r (net181),
    .q (net190),
    .notq (net189)
  );
  and_cell and52 (
    .a (net182),
    .b (net184),
    .out (net191)
  );
  and_cell and53 (
    .a (net191),
    .b (net186),
    .out (net192)
  );
  and_cell and54 (
    .a (net192),
    .b (net188),
    .out (net193)
  );
  and_cell and55 (
    .a (net193),
    .b (net190),
    .out (net194)
  );
  dffsr_cell flop71 (
    .d (net196),
    .clk (net146),
    .s (net197),
    .r (net197),
    .q (net198),
    .notq (net196)
  );
  dffsr_cell flop72 (
    .d (net199),
    .clk (net196),
    .s (net197),
    .r (net197),
    .q (net200),
    .notq (net199)
  );
  dffsr_cell flop73 (
    .d (net201),
    .clk (net199),
    .s (net197),
    .r (net197),
    .q (net202),
    .notq (net201)
  );
  dffsr_cell flop74 (
    .d (net203),
    .clk (net201),
    .s (net197),
    .r (net197),
    .q (net204),
    .notq (net203)
  );
  dffsr_cell flop75 (
    .d (net205),
    .clk (net203),
    .s (net197),
    .r (net197),
    .q (net206),
    .notq (net205)
  );
  and_cell and56 (
    .a (net198),
    .b (net200),
    .out (net207)
  );
  and_cell and57 (
    .a (net207),
    .b (net202),
    .out (net208)
  );
  and_cell and58 (
    .a (net208),
    .b (net204),
    .out (net209)
  );
  and_cell and59 (
    .a (net209),
    .b (net206),
    .out (net210)
  );
  dffsr_cell flop76 (
    .d (net212),
    .clk (net162),
    .s (net213),
    .r (net213),
    .q (net214),
    .notq (net212)
  );
  dffsr_cell flop77 (
    .d (net215),
    .clk (net212),
    .s (net213),
    .r (net213),
    .q (net216),
    .notq (net215)
  );
  dffsr_cell flop78 (
    .d (net217),
    .clk (net215),
    .s (net213),
    .r (net213),
    .q (net218),
    .notq (net217)
  );
  dffsr_cell flop79 (
    .d (net219),
    .clk (net217),
    .s (net213),
    .r (net213),
    .q (net220),
    .notq (net219)
  );
  dffsr_cell flop80 (
    .d (net221),
    .clk (net219),
    .s (net213),
    .r (net213),
    .q (net222),
    .notq (net221)
  );
  and_cell and60 (
    .a (net214),
    .b (net216),
    .out (net223)
  );
  and_cell and61 (
    .a (net223),
    .b (net218),
    .out (net224)
  );
  and_cell and62 (
    .a (net224),
    .b (net220),
    .out (net225)
  );
  and_cell and63 (
    .a (net225),
    .b (net222),
    .out (net226)
  );
  dffsr_cell flop81 (
    .d (net228),
    .clk (net1),
    .s (net229),
    .r (net229),
    .q (net230),
    .notq (net228)
  );
  dffsr_cell flop82 (
    .d (net231),
    .clk (net228),
    .s (net229),
    .r (net229),
    .q (net232),
    .notq (net231)
  );
  dffsr_cell flop83 (
    .d (net233),
    .clk (net231),
    .s (net229),
    .r (net229),
    .q (net234),
    .notq (net233)
  );
  dffsr_cell flop84 (
    .d (net235),
    .clk (net233),
    .s (net229),
    .r (net229),
    .q (net236),
    .notq (net235)
  );
  dffsr_cell flop85 (
    .d (net237),
    .clk (net235),
    .s (net229),
    .r (net229),
    .q (net238),
    .notq (net237)
  );
  and_cell and64 (
    .a (net230),
    .b (net232),
    .out (net239)
  );
  and_cell and65 (
    .a (net239),
    .b (net234),
    .out (net240)
  );
  and_cell and66 (
    .a (net240),
    .b (net236),
    .out (net241)
  );
  and_cell and67 (
    .a (net241),
    .b (net238),
    .out (net242)
  );
  dffsr_cell flop86 (
    .d (net244),
    .clk (net242),
    .s (net245),
    .r (net245),
    .q (net246),
    .notq (net244)
  );
  dffsr_cell flop87 (
    .d (net247),
    .clk (net244),
    .s (net245),
    .r (net245),
    .q (net248),
    .notq (net247)
  );
  dffsr_cell flop88 (
    .d (net249),
    .clk (net247),
    .s (net245),
    .r (net245),
    .q (net250),
    .notq (net249)
  );
  dffsr_cell flop89 (
    .d (net251),
    .clk (net249),
    .s (net245),
    .r (net245),
    .q (net252),
    .notq (net251)
  );
  dffsr_cell flop90 (
    .d (net253),
    .clk (net251),
    .s (net245),
    .r (net245),
    .q (net254),
    .notq (net253)
  );
  and_cell and68 (
    .a (net246),
    .b (net248),
    .out (net255)
  );
  and_cell and69 (
    .a (net255),
    .b (net250),
    .out (net256)
  );
  and_cell and70 (
    .a (net256),
    .b (net252),
    .out (net257)
  );
  and_cell and71 (
    .a (net257),
    .b (net254),
    .out (net258)
  );
  mux_cell mux1 (
    .a (net1),
    .b (net3),
    .sel (net4),
    .out (net16)
  );
  or_cell or1 (
    .a (net178),
    .b (net194),
    .out (net261)
  );
  or_cell or2 (
    .a (net261),
    .b (net210),
    .out (net262)
  );
  or_cell or3 (
    .a (net262),
    .b (net226),
    .out (net263)
  );
  or_cell or4 (
    .a (net263),
    .b (net258),
    .out (net19)
  );
  dffsr_cell flop91 (
    .d (net264),
    .clk (net1),
    .s (net265),
    .r (net265),
    .q (net266),
    .notq (net264)
  );
  dffsr_cell flop92 (
    .d (net267),
    .clk (net264),
    .s (net265),
    .r (net265),
    .q (net268),
    .notq (net267)
  );
  and_cell and73 (
    .a (net266),
    .b (net268),
    .out (net269)
  );
  dffsr_cell flop93 (
    .d (net271),
    .clk (net269),
    .s (net272),
    .r (net272),
    .q (net273),
    .notq (net271)
  );
  dffsr_cell flop94 (
    .d (net274),
    .clk (net271),
    .s (net272),
    .r (net272),
    .q (net275),
    .notq (net274)
  );
  and_cell and74 (
    .a (net273),
    .b (net275),
    .out (net276)
  );
  dffsr_cell flop95 (
    .d (net278),
    .clk (net269),
    .s (net279),
    .r (net279),
    .q (net280),
    .notq (net278)
  );
  dffsr_cell flop96 (
    .d (net281),
    .clk (net278),
    .s (net279),
    .r (net279),
    .q (net282),
    .notq (net281)
  );
  and_cell and72 (
    .a (net280),
    .b (net282),
    .out (net283)
  );
  dffsr_cell flop97 (
    .d (net285),
    .clk (net269),
    .s (net286),
    .r (net286),
    .q (net287),
    .notq (net285)
  );
  dffsr_cell flop98 (
    .d (net288),
    .clk (net285),
    .s (net286),
    .r (net286),
    .q (net289),
    .notq (net288)
  );
  and_cell and75 (
    .a (net287),
    .b (net289),
    .out (net290)
  );
  dffsr_cell flop99 (
    .d (net292),
    .clk (net276),
    .s (net293),
    .r (net293),
    .q (net294),
    .notq (net292)
  );
  dffsr_cell flop100 (
    .d (net295),
    .clk (net292),
    .s (net293),
    .r (net293),
    .q (net296),
    .notq (net295)
  );
  and_cell and76 (
    .a (net294),
    .b (net296),
    .out (net297)
  );
  dffsr_cell flop101 (
    .d (net299),
    .clk (net290),
    .s (net300),
    .r (net300),
    .q (net301),
    .notq (net299)
  );
  dffsr_cell flop102 (
    .d (net302),
    .clk (net299),
    .s (net300),
    .r (net300),
    .q (net303),
    .notq (net302)
  );
  dffsr_cell flop103 (
    .d (net304),
    .clk (net302),
    .s (net300),
    .r (net300),
    .q (net305),
    .notq (net304)
  );
  and_cell and77 (
    .a (net301),
    .b (net303),
    .out (net306)
  );
  and_cell and78 (
    .a (net306),
    .b (net305),
    .out (net307)
  );
  dffsr_cell flop104 (
    .d (net309),
    .clk (net283),
    .s (net310),
    .r (net310),
    .q (net311),
    .notq (net309)
  );
  dffsr_cell flop105 (
    .d (net312),
    .clk (net309),
    .s (net310),
    .r (net310),
    .q (net313),
    .notq (net312)
  );
  and_cell and79 (
    .a (net311),
    .b (net313),
    .out (net314)
  );
  or_cell or5 (
    .a (net297),
    .b (net307),
    .out (net316)
  );
  or_cell or6 (
    .a (net316),
    .b (net314),
    .out (net31)
  );
  dffsr_cell flop5 (
    .d (net317),
    .clk (net9),
    .s (net318),
    .r (net318),
    .q (net319),
    .notq (net317)
  );
  dffsr_cell flop6 (
    .d (net320),
    .clk (net317),
    .s (net318),
    .r (net318),
    .q (net321),
    .notq (net320)
  );
  and_cell and1 (
    .a (net319),
    .b (net321),
    .out (net322)
  );
  dffsr_cell flop7 (
    .d (net324),
    .clk (net8),
    .s (net325),
    .r (net325),
    .q (net326),
    .notq (net324)
  );
  dffsr_cell flop8 (
    .d (net327),
    .clk (net324),
    .s (net325),
    .r (net325),
    .q (net328),
    .notq (net327)
  );
  dffsr_cell flop9 (
    .d (net329),
    .clk (net327),
    .s (net325),
    .r (net325),
    .q (net330),
    .notq (net329)
  );
  and_cell and3 (
    .a (net326),
    .b (net328),
    .out (net331)
  );
  and_cell and5 (
    .a (net331),
    .b (net330),
    .out (net332)
  );
  dffsr_cell flop10 (
    .d (net335),
    .clk (net7),
    .s (net336),
    .r (net336),
    .q (net337),
    .notq (net335)
  );
  dffsr_cell flop11 (
    .d (net338),
    .clk (net335),
    .s (net336),
    .r (net336),
    .q (net339),
    .notq (net338)
  );
  and_cell and6 (
    .a (net337),
    .b (net339),
    .out (net340)
  );
  dffsr_cell flop12 (
    .d (net342),
    .clk (net6),
    .s (net343),
    .r (net343),
    .q (net344),
    .notq (net342)
  );
  dffsr_cell flop13 (
    .d (net345),
    .clk (net342),
    .s (net343),
    .r (net343),
    .q (net346),
    .notq (net345)
  );
  dffsr_cell flop14 (
    .d (net347),
    .clk (net345),
    .s (net343),
    .r (net343),
    .q (net348),
    .notq (net347)
  );
  and_cell and7 (
    .a (net344),
    .b (net346),
    .out (net349)
  );
  and_cell and8 (
    .a (net349),
    .b (net348),
    .out (net350)
  );
  dffsr_cell flop15 (
    .d (net352),
    .clk (net322),
    .s (net353),
    .r (net353),
    .q (net354),
    .notq (net352)
  );
  dffsr_cell flop36 (
    .d (net355),
    .clk (net352),
    .s (net353),
    .r (net353),
    .q (net356),
    .notq (net355)
  );
  and_cell and9 (
    .a (net354),
    .b (net356),
    .out (net357)
  );
  dffsr_cell flop37 (
    .d (net359),
    .clk (net332),
    .s (net360),
    .r (net360),
    .q (net361),
    .notq (net359)
  );
  dffsr_cell flop38 (
    .d (net362),
    .clk (net359),
    .s (net360),
    .r (net360),
    .q (net363),
    .notq (net362)
  );
  dffsr_cell flop39 (
    .d (net364),
    .clk (net362),
    .s (net360),
    .r (net360),
    .q (net365),
    .notq (net364)
  );
  and_cell and26 (
    .a (net361),
    .b (net363),
    .out (net366)
  );
  and_cell and27 (
    .a (net366),
    .b (net365),
    .out (net367)
  );
  dffsr_cell flop106 (
    .d (net369),
    .clk (net340),
    .s (net370),
    .r (net370),
    .q (net371),
    .notq (net369)
  );
  dffsr_cell flop107 (
    .d (net372),
    .clk (net369),
    .s (net370),
    .r (net370),
    .q (net373),
    .notq (net372)
  );
  and_cell and28 (
    .a (net371),
    .b (net373),
    .out (net374)
  );
  dffsr_cell flop108 (
    .d (net376),
    .clk (net350),
    .s (net377),
    .r (net377),
    .q (net378),
    .notq (net376)
  );
  dffsr_cell flop109 (
    .d (net379),
    .clk (net376),
    .s (net377),
    .r (net377),
    .q (net380),
    .notq (net379)
  );
  dffsr_cell flop110 (
    .d (net381),
    .clk (net379),
    .s (net377),
    .r (net377),
    .q (net382),
    .notq (net381)
  );
  and_cell and29 (
    .a (net378),
    .b (net380),
    .out (net383)
  );
  and_cell and30 (
    .a (net383),
    .b (net382),
    .out (net384)
  );
  dffsr_cell flop111 (
    .d (net386),
    .clk (net387),
    .s (net388),
    .r (net388),
    .q (net389),
    .notq (net386)
  );
  dffsr_cell flop112 (
    .d (net390),
    .clk (net386),
    .s (net388),
    .r (net388),
    .q (net391),
    .notq (net390)
  );
  dffsr_cell flop113 (
    .d (net392),
    .clk (net390),
    .s (net388),
    .r (net388),
    .q (net393),
    .notq (net392)
  );
  dffsr_cell flop114 (
    .d (net394),
    .clk (net392),
    .s (net388),
    .r (net388),
    .q (net395),
    .notq (net394)
  );
  dffsr_cell flop115 (
    .d (net396),
    .clk (net394),
    .s (net388),
    .r (net388),
    .q (net397),
    .notq (net396)
  );
  dffsr_cell flop116 (
    .d (net398),
    .clk (net396),
    .s (net388),
    .r (net388),
    .q (net399),
    .notq (net398)
  );
  and_cell and31 (
    .a (net389),
    .b (net391),
    .out (net400)
  );
  and_cell and32 (
    .a (net400),
    .b (net393),
    .out (net401)
  );
  and_cell and33 (
    .a (net401),
    .b (net402),
    .out (net403)
  );
  and_cell and34 (
    .a (net395),
    .b (net397),
    .out (net404)
  );
  and_cell and80 (
    .a (net404),
    .b (net399),
    .out (net402)
  );
  dffsr_cell flop117 (
    .d (net405),
    .clk (net406),
    .s (net407),
    .r (net407),
    .q (net408),
    .notq (net405)
  );
  dffsr_cell flop118 (
    .d (net409),
    .clk (net405),
    .s (net407),
    .r (net407),
    .q (net410),
    .notq (net409)
  );
  dffsr_cell flop119 (
    .d (net411),
    .clk (net409),
    .s (net407),
    .r (net407),
    .q (net412),
    .notq (net411)
  );
  dffsr_cell flop120 (
    .d (net413),
    .clk (net411),
    .s (net407),
    .r (net407),
    .q (net414),
    .notq (net413)
  );
  dffsr_cell flop121 (
    .d (net415),
    .clk (net413),
    .s (net407),
    .r (net407),
    .q (net416),
    .notq (net415)
  );
  and_cell and81 (
    .a (net408),
    .b (net410),
    .out (net417)
  );
  and_cell and82 (
    .a (net417),
    .b (net412),
    .out (net418)
  );
  and_cell and83 (
    .a (net418),
    .b (net414),
    .out (net419)
  );
  and_cell and84 (
    .a (net419),
    .b (net416),
    .out (net420)
  );
  dffsr_cell flop122 (
    .d (net422),
    .clk (net374),
    .s (net423),
    .r (net423),
    .q (net424),
    .notq (net422)
  );
  dffsr_cell flop123 (
    .d (net425),
    .clk (net422),
    .s (net423),
    .r (net423),
    .q (net426),
    .notq (net425)
  );
  dffsr_cell flop124 (
    .d (net427),
    .clk (net425),
    .s (net423),
    .r (net423),
    .q (net428),
    .notq (net427)
  );
  and_cell and85 (
    .a (net424),
    .b (net426),
    .out (net429)
  );
  and_cell and86 (
    .a (net429),
    .b (net428),
    .out (net430)
  );
  dffsr_cell flop125 (
    .d (net432),
    .clk (net384),
    .s (net433),
    .r (net433),
    .q (net434),
    .notq (net432)
  );
  dffsr_cell flop126 (
    .d (net435),
    .clk (net432),
    .s (net433),
    .r (net433),
    .q (net436),
    .notq (net435)
  );
  dffsr_cell flop127 (
    .d (net437),
    .clk (net435),
    .s (net433),
    .r (net433),
    .q (net438),
    .notq (net437)
  );
  dffsr_cell flop128 (
    .d (net439),
    .clk (net437),
    .s (net433),
    .r (net433),
    .q (net440),
    .notq (net439)
  );
  dffsr_cell flop129 (
    .d (net441),
    .clk (net439),
    .s (net433),
    .r (net433),
    .q (net442),
    .notq (net441)
  );
  and_cell and87 (
    .a (net434),
    .b (net436),
    .out (net443)
  );
  and_cell and88 (
    .a (net443),
    .b (net438),
    .out (net444)
  );
  and_cell and89 (
    .a (net444),
    .b (net440),
    .out (net445)
  );
  and_cell and90 (
    .a (net445),
    .b (net442),
    .out (net446)
  );
  dffsr_cell flop130 (
    .d (net448),
    .clk (net420),
    .s (net449),
    .r (net449),
    .q (net450),
    .notq (net448)
  );
  dffsr_cell flop131 (
    .d (net451),
    .clk (net448),
    .s (net449),
    .r (net449),
    .q (net452),
    .notq (net451)
  );
  dffsr_cell flop132 (
    .d (net453),
    .clk (net451),
    .s (net449),
    .r (net449),
    .q (net454),
    .notq (net453)
  );
  and_cell and91 (
    .a (net450),
    .b (net452),
    .out (net455)
  );
  and_cell and92 (
    .a (net455),
    .b (net454),
    .out (net456)
  );
  dffsr_cell flop133 (
    .d (net458),
    .clk (net403),
    .s (net459),
    .r (net459),
    .q (net460),
    .notq (net458)
  );
  dffsr_cell flop134 (
    .d (net461),
    .clk (net458),
    .s (net459),
    .r (net459),
    .q (net462),
    .notq (net461)
  );
  dffsr_cell flop135 (
    .d (net463),
    .clk (net461),
    .s (net459),
    .r (net459),
    .q (net464),
    .notq (net463)
  );
  dffsr_cell flop136 (
    .d (net465),
    .clk (net463),
    .s (net459),
    .r (net459),
    .q (net466),
    .notq (net465)
  );
  dffsr_cell flop137 (
    .d (net467),
    .clk (net465),
    .s (net459),
    .r (net459),
    .q (net468),
    .notq (net467)
  );
  and_cell and93 (
    .a (net460),
    .b (net462),
    .out (net469)
  );
  and_cell and94 (
    .a (net469),
    .b (net464),
    .out (net470)
  );
  and_cell and95 (
    .a (net470),
    .b (net466),
    .out (net471)
  );
  and_cell and96 (
    .a (net471),
    .b (net468),
    .out (net472)
  );
  dffsr_cell flop138 (
    .d (net474),
    .clk (net357),
    .s (net475),
    .r (net475),
    .q (net476),
    .notq (net474)
  );
  dffsr_cell flop139 (
    .d (net477),
    .clk (net474),
    .s (net475),
    .r (net475),
    .q (net478),
    .notq (net477)
  );
  dffsr_cell flop140 (
    .d (net479),
    .clk (net477),
    .s (net475),
    .r (net475),
    .q (net480),
    .notq (net479)
  );
  and_cell and97 (
    .a (net476),
    .b (net478),
    .out (net481)
  );
  and_cell and98 (
    .a (net481),
    .b (net480),
    .out (net482)
  );
  dffsr_cell flop141 (
    .d (net484),
    .clk (net367),
    .s (net485),
    .r (net485),
    .q (net486),
    .notq (net484)
  );
  dffsr_cell flop142 (
    .d (net487),
    .clk (net484),
    .s (net485),
    .r (net485),
    .q (net488),
    .notq (net487)
  );
  dffsr_cell flop143 (
    .d (net489),
    .clk (net487),
    .s (net485),
    .r (net485),
    .q (net490),
    .notq (net489)
  );
  dffsr_cell flop144 (
    .d (net491),
    .clk (net489),
    .s (net485),
    .r (net485),
    .q (net492),
    .notq (net491)
  );
  dffsr_cell flop145 (
    .d (net493),
    .clk (net491),
    .s (net485),
    .r (net485),
    .q (net494),
    .notq (net493)
  );
  and_cell and99 (
    .a (net486),
    .b (net488),
    .out (net495)
  );
  and_cell and100 (
    .a (net495),
    .b (net490),
    .out (net496)
  );
  and_cell and101 (
    .a (net496),
    .b (net492),
    .out (net497)
  );
  and_cell and102 (
    .a (net497),
    .b (net494),
    .out (net498)
  );
  dffsr_cell flop146 (
    .d (net500),
    .clk (net27),
    .s (net501),
    .r (net501),
    .q (net502),
    .notq (net500)
  );
  dffsr_cell flop147 (
    .d (net503),
    .clk (net500),
    .s (net501),
    .r (net501),
    .q (net504),
    .notq (net503)
  );
  and_cell and106 (
    .a (net502),
    .b (net504),
    .out (net406)
  );
  dffsr_cell flop148 (
    .d (net506),
    .clk (net29),
    .s (net507),
    .r (net507),
    .q (net508),
    .notq (net506)
  );
  dffsr_cell flop149 (
    .d (net509),
    .clk (net506),
    .s (net507),
    .r (net507),
    .q (net510),
    .notq (net509)
  );
  dffsr_cell flop150 (
    .d (net511),
    .clk (net509),
    .s (net507),
    .r (net507),
    .q (net512),
    .notq (net511)
  );
  and_cell and107 (
    .a (net508),
    .b (net510),
    .out (net513)
  );
  and_cell and108 (
    .a (net513),
    .b (net512),
    .out (net387)
  );
  or_cell or7 (
    .a (net482),
    .b (net498),
    .out (net21)
  );
  or_cell or8 (
    .a (net430),
    .b (net446),
    .out (net23)
  );
  or_cell or9 (
    .a (net456),
    .b (net472),
    .out (net516)
  );
  dffsr_cell flop151 (
    .d (net517),
    .clk (net16),
    .s (net518),
    .r (net518),
    .q (net519),
    .notq (net517)
  );
  dffsr_cell flop152 (
    .d (net520),
    .clk (net517),
    .s (net518),
    .r (net518),
    .q (net521),
    .notq (net520)
  );
  dffsr_cell flop153 (
    .d (net522),
    .clk (net520),
    .s (net518),
    .r (net518),
    .q (net523),
    .notq (net522)
  );
  and_cell and103 (
    .a (net519),
    .b (net521),
    .out (net524)
  );
  and_cell and104 (
    .a (net524),
    .b (net523),
    .out (net525)
  );
  dffsr_cell flop154 (
    .d (net527),
    .clk (net528),
    .s (net529),
    .r (net529),
    .q (net530),
    .notq (net527)
  );
  dffsr_cell flop155 (
    .d (net531),
    .clk (net527),
    .s (net529),
    .r (net529),
    .q (net532),
    .notq (net531)
  );
  dffsr_cell flop156 (
    .d (net533),
    .clk (net531),
    .s (net529),
    .r (net529),
    .q (net534),
    .notq (net533)
  );
  and_cell and105 (
    .a (net530),
    .b (net532),
    .out (net535)
  );
  and_cell and109 (
    .a (net535),
    .b (net534),
    .out (net536)
  );
  dffsr_cell flop157 (
    .d (net528),
    .clk (net525),
    .s (net538),
    .r (net538),
    .q (net539),
    .notq (net528)
  );
  dffsr_cell flop158 (
    .d (net540),
    .clk (net528),
    .s (net538),
    .r (net538),
    .q (net541),
    .notq (net540)
  );
  dffsr_cell flop159 (
    .d (net542),
    .clk (net540),
    .s (net538),
    .r (net538),
    .q (net543),
    .notq (net542)
  );
  and_cell and110 (
    .a (net539),
    .b (net541),
    .out (net544)
  );
  and_cell and111 (
    .a (net544),
    .b (net543),
    .out (net545)
  );
  dffsr_cell flop160 (
    .d (net547),
    .clk (net525),
    .s (net548),
    .r (net548),
    .q (net549),
    .notq (net547)
  );
  dffsr_cell flop161 (
    .d (net550),
    .clk (net547),
    .s (net548),
    .r (net548),
    .q (net551),
    .notq (net550)
  );
  dffsr_cell flop162 (
    .d (net552),
    .clk (net550),
    .s (net548),
    .r (net548),
    .q (net553),
    .notq (net552)
  );
  and_cell and112 (
    .a (net549),
    .b (net551),
    .out (net554)
  );
  and_cell and113 (
    .a (net554),
    .b (net553),
    .out (net555)
  );
  dffsr_cell flop163 (
    .d (net557),
    .clk (net536),
    .s (net558),
    .r (net558),
    .q (net559),
    .notq (net557)
  );
  dffsr_cell flop164 (
    .d (net560),
    .clk (net557),
    .s (net558),
    .r (net558),
    .q (net561),
    .notq (net560)
  );
  dffsr_cell flop165 (
    .d (net562),
    .clk (net560),
    .s (net558),
    .r (net558),
    .q (net563),
    .notq (net562)
  );
  and_cell and114 (
    .a (net559),
    .b (net561),
    .out (net564)
  );
  and_cell and115 (
    .a (net564),
    .b (net563),
    .out (net565)
  );
  dffsr_cell flop166 (
    .d (net567),
    .clk (net568),
    .s (net569),
    .r (net569),
    .q (net570),
    .notq (net567)
  );
  dffsr_cell flop167 (
    .d (net571),
    .clk (net567),
    .s (net569),
    .r (net569),
    .q (net572),
    .notq (net571)
  );
  dffsr_cell flop168 (
    .d (net573),
    .clk (net571),
    .s (net569),
    .r (net569),
    .q (net574),
    .notq (net573)
  );
  and_cell and116 (
    .a (net570),
    .b (net572),
    .out (net575)
  );
  and_cell and117 (
    .a (net575),
    .b (net574),
    .out (net576)
  );
  dffsr_cell flop169 (
    .d (net578),
    .clk (net579),
    .s (net580),
    .r (net580),
    .q (net581),
    .notq (net578)
  );
  dffsr_cell flop170 (
    .d (net582),
    .clk (net578),
    .s (net580),
    .r (net580),
    .q (net583),
    .notq (net582)
  );
  dffsr_cell flop171 (
    .d (net584),
    .clk (net582),
    .s (net580),
    .r (net580),
    .q (net585),
    .notq (net584)
  );
  and_cell and118 (
    .a (net581),
    .b (net583),
    .out (net586)
  );
  and_cell and119 (
    .a (net586),
    .b (net585),
    .out (net587)
  );
  or_cell or10 (
    .a (net545),
    .b (net555),
    .out (net568)
  );
  or_cell or11 (
    .a (net565),
    .b (net576),
    .out (net579)
  );
  mux_cell mux2 (
    .a (net516),
    .b (net587),
    .sel (net5),
    .out (net25)
  );
endmodule
