/* Automatically generated from https://wokwi.com/projects/377426511818305537 */

`default_nettype none

module tt_um_wokwi_377426511818305537(
  input  wire [7:0] ui_in,    // Dedicated inputs
  output wire [7:0] uo_out,    // Dedicated outputs
  input  wire [7:0] uio_in,    // IOs: Input path
  output wire [7:0] uio_out,    // IOs: Output path
  output wire [7:0] uio_oe,    // IOs: Enable path (active high: 0=input, 1=output)
  input ena,
  input clk,
  input rst_n
);
  wire net1 = clk;
  wire net2 = rst_n;
  wire net3 = ui_in[0];
  wire net4 = ui_in[1];
  wire net5 = ui_in[2];
  wire net6 = ui_in[3];
  wire net7 = ui_in[4];
  wire net8 = ui_in[7];
  wire net9;
  wire net10;
  wire net11;
  wire net12;
  wire net13;
  wire net14;
  wire net15;
  wire net16;
  wire net17;
  wire net18 = 1'b1;
  wire net19;
  wire net20;
  wire net21;
  wire net22;
  wire net23;
  wire net24;
  wire net25;
  wire net26;
  wire net27;
  wire net28;
  wire net29;
  wire net30;
  wire net31;
  wire net32;
  wire net33;
  wire net34;
  wire net35;
  wire net36;
  wire net37;
  wire net38;
  wire net39;
  wire net40;
  wire net41;
  wire net42;
  wire net43;
  wire net44;
  wire net45;
  wire net46;
  wire net47;
  wire net48;
  wire net49;
  wire net50;
  wire net51;
  wire net52;
  wire net53;
  wire net54;
  wire net55;
  wire net56;
  wire net57;
  wire net58;
  wire net59;
  wire net60;
  wire net61;
  wire net62;
  wire net63;
  wire net64;
  wire net65;
  wire net66;
  wire net67;
  wire net68;
  wire net69;
  wire net70;
  wire net71;
  wire net72;
  wire net73;
  wire net74;
  wire net75;
  wire net76;
  wire net77;
  wire net78;
  wire net79;
  wire net80;
  wire net81;
  wire net82;
  wire net83 = 1'b1;
  wire net84 = 1'b1;
  wire net85 = 1'b0;
  wire net86 = 1'b1;
  wire net87 = 1'b0;
  wire net88;
  wire net89;
  wire net90;
  wire net91;
  wire net92;
  wire net93;
  wire net94;
  wire net95;
  wire net96;
  wire net97;
  wire net98;
  wire net99;
  wire net100 = 1'b0;
  wire net101;
  wire net102;
  wire net103;
  wire net104;
  wire net105;
  wire net106;
  wire net107;
  wire net108;
  wire net109;
  wire net110;
  wire net111;
  wire net112;
  wire net113;
  wire net114;
  wire net115;
  wire net116;
  wire net117 = 1'b0;
  wire net118;
  wire net119;
  wire net120;
  wire net121;
  wire net122;
  wire net123;
  wire net124;
  wire net125;
  wire net126;
  wire net127;
  wire net128;
  wire net129;
  wire net130;
  wire net131;
  wire net132;
  wire net133;
  wire net134;
  wire net135;
  wire net136;
  wire net137;
  wire net138;
  wire net139;
  wire net140;
  wire net141;
  wire net142;
  wire net143;
  wire net144;
  wire net145;
  wire net146;
  wire net147;
  wire net148;
  wire net149;
  wire net150;
  wire net151;
  wire net152;
  wire net153;
  wire net154;
  wire net155;
  wire net156;
  wire net157;
  wire net158;
  wire net159;
  wire net160;
  wire net161;
  wire net162;
  wire net163;
  wire net164;
  wire net165;
  wire net166;
  wire net167;
  wire net168;
  wire net169;
  wire net170;
  wire net171;
  wire net172;
  wire net173;
  wire net174;
  wire net175 = 1'b0;
  wire net176;
  wire net177;
  wire net178 = 1'b0;
  wire net179;
  wire net180;
  wire net181;
  wire net182;
  wire net183;
  wire net184;
  wire net185;
  wire net186;
  wire net187;
  wire net188;
  wire net189;
  wire net190;
  wire net191;
  wire net192;
  wire net193;
  wire net194;
  wire net195;
  wire net196;
  wire net197;
  wire net198;
  wire net199;
  wire net200;
  wire net201;
  wire net202;
  wire net203;
  wire net204;
  wire net205;
  wire net206;
  wire net207;
  wire net208;
  wire net209;
  wire net210;
  wire net211;
  wire net212;
  wire net213;
  wire net214;
  wire net215;
  wire net216;
  wire net217;
  wire net218;
  wire net219;
  wire net220;
  wire net221;
  wire net222;
  wire net223;
  wire net224;
  wire net225;
  wire net226;
  wire net227;
  wire net228;
  wire net229;
  wire net230;
  wire net231;
  wire net232;
  wire net233;
  wire net234;
  wire net235;
  wire net236;
  wire net237;
  wire net238;
  wire net239;
  wire net240;
  wire net241;
  wire net242;
  wire net243;
  wire net244;
  wire net245;
  wire net246;
  wire net247;
  wire net248;
  wire net249;
  wire net250;
  wire net251;
  wire net252 = 1'b0;
  wire net253;
  wire net254;
  wire net255;
  wire net256 = 1'b0;
  wire net257;
  wire net258;
  wire net259;
  wire net260;
  wire net261;
  wire net262;
  wire net263;
  wire net264;
  wire net265;
  wire net266;
  wire net267;
  wire net268;
  wire net269;
  wire net270;
  wire net271;
  wire net272;
  wire net273;
  wire net274;
  wire net275;
  wire net276;
  wire net277;
  wire net278;
  wire net279;
  wire net280;
  wire net281;
  wire net282;
  wire net283;
  wire net284;
  wire net285;
  wire net286;
  wire net287;
  wire net288;
  wire net289;
  wire net290;
  wire net291;
  wire net292;
  wire net293;
  wire net294;
  wire net295;
  wire net296;
  wire net297;
  wire net298;
  wire net299;
  wire net300;
  wire net301;
  wire net302;
  wire net303;
  wire net304;
  wire net305;
  wire net306;
  wire net307;
  wire net308;
  wire net309;
  wire net310;
  wire net311;
  wire net312;
  wire net313;
  wire net314;
  wire net315;
  wire net316;
  wire net317;
  wire net318;
  wire net319;
  wire net320;
  wire net321;
  wire net322;
  wire net323;
  wire net324;
  wire net325;
  wire net326;
  wire net327;
  wire net328;
  wire net329;
  wire net330 = 1'b0;
  wire net331;
  wire net332;
  wire net333 = 1'b0;
  wire net334;
  wire net335;
  wire net336 = 1'b0;
  wire net337;
  wire net338 = 1'b1;
  wire net339;
  wire net340 = 1'b0;
  wire net341 = 1'b0;
  wire net342 = 1'b0;
  wire net343;
  wire net344;
  wire net345;
  wire net346;
  wire net347;
  wire net348;
  wire net349;
  wire net350;
  wire net351;
  wire net352;
  wire net353;
  wire net354;
  wire net355;
  wire net356;
  wire net357;
  wire net358;
  wire net359;
  wire net360;
  wire net361;
  wire net362;
  wire net363;
  wire net364;
  wire net365;
  wire net366;

  assign uo_out[0] = net9;
  assign uo_out[1] = net10;
  assign uo_out[2] = net11;
  assign uo_out[3] = net12;
  assign uo_out[4] = net13;
  assign uo_out[5] = net14;
  assign uo_out[6] = net15;
  assign uo_out[7] = net16;
  assign uio_out[0] = net17;
  assign uio_oe[0] = net18;
  assign uio_out[1] = net19;
  assign uio_oe[1] = net18;
  assign uio_out[2] = net20;
  assign uio_oe[2] = net18;
  assign uio_out[3] = net21;
  assign uio_oe[3] = net18;
  assign uio_out[4] = net13;
  assign uio_oe[4] = net18;
  assign uio_out[5] = net22;
  assign uio_oe[5] = net18;
  assign uio_out[6] = net23;
  assign uio_oe[6] = net18;
  assign uio_out[7] = 0;
  assign uio_oe[7] = net18;

  mux_cell mux1 (
    .a (net24),
    .b (net25),
    .sel (net26),
    .out (net27)
  );
  mux_cell mux2 (
    .a (net28),
    .b (net29),
    .sel (net30),
    .out (net24)
  );
  xor_cell xor1 (
    .a (net29),
    .b (net31),
    .out (net25)
  );
  mux_cell mux3 (
    .a (net32),
    .b (net33),
    .sel (net34),
    .out (net35)
  );
  mux_cell mux4 (
    .a (net36),
    .b (net37),
    .sel (net38),
    .out (net39)
  );
  mux_cell mux5 (
    .a (net27),
    .b (net40),
    .sel (net41),
    .out (net32)
  );
  mux_cell mux6 (
    .a (net35),
    .b (net42),
    .sel (net43),
    .out (net36)
  );
  xor_cell xor2 (
    .a (net40),
    .b (net31),
    .out (net33)
  );
  xor_cell xor3 (
    .a (net42),
    .b (net31),
    .out (net37)
  );
  mux_cell mux7 (
    .a (net44),
    .b (net45),
    .sel (net46),
    .out (net47)
  );
  mux_cell mux8 (
    .a (net48),
    .b (net49),
    .sel (net50),
    .out (net51)
  );
  mux_cell mux9 (
    .a (net52),
    .b (net53),
    .sel (net54),
    .out (net55)
  );
  mux_cell mux10 (
    .a (net56),
    .b (net57),
    .sel (net58),
    .out (net59)
  );
  mux_cell mux11 (
    .a (net39),
    .b (net60),
    .sel (net61),
    .out (net44)
  );
  mux_cell mux12 (
    .a (net47),
    .b (net62),
    .sel (net63),
    .out (net48)
  );
  mux_cell mux13 (
    .a (net51),
    .b (net64),
    .sel (net65),
    .out (net52)
  );
  mux_cell mux14 (
    .a (net55),
    .b (net66),
    .sel (net67),
    .out (net56)
  );
  xor_cell xor4 (
    .a (net60),
    .b (net31),
    .out (net45)
  );
  xor_cell xor5 (
    .a (net62),
    .b (net31),
    .out (net49)
  );
  xor_cell xor6 (
    .a (net64),
    .b (net31),
    .out (net53)
  );
  xor_cell xor7 (
    .a (net66),
    .b (net31),
    .out (net57)
  );
  and_cell and1 (
    .a (net31),
    .b (net68),
    .out (net69)
  );
  and_cell and2 (
    .a (net69),
    .b (net70),
    .out (net71)
  );
  and_cell and3 (
    .a (net71),
    .b (net72),
    .out (net73)
  );
  and_cell and4 (
    .a (net73),
    .b (net74),
    .out (net75)
  );
  and_cell and5 (
    .a (net75),
    .b (net76),
    .out (net77)
  );
  and_cell and6 (
    .a (net77),
    .b (net78),
    .out (net79)
  );
  and_cell and7 (
    .a (net79),
    .b (net80),
    .out (net81)
  );
  or_cell or1 (
    .a (net81),
    .b (net31),
    .out (net28)
  );
  not_cell not1 (
    .in (net2),
    .out (net82)
  );
  and_cell and8 (
    .a (net67),
    .b (net88),
    .out (net58)
  );
  and_cell and9 (
    .a (net65),
    .b (net89),
    .out (net54)
  );
  and_cell and10 (
    .a (net63),
    .b (net90),
    .out (net50)
  );
  and_cell and11 (
    .a (net61),
    .b (net91),
    .out (net46)
  );
  and_cell and12 (
    .a (net43),
    .b (net92),
    .out (net38)
  );
  and_cell and13 (
    .a (net41),
    .b (net93),
    .out (net34)
  );
  and_cell and14 (
    .a (net30),
    .b (net94),
    .out (net26)
  );
  dffsr_cell flop1 (
    .d (net95),
    .clk (net96),
    .s (net8),
    .r (net82),
    .q (net97)
  );
  dffsr_cell flop2 (
    .d (net97),
    .clk (net96),
    .s (net8),
    .r (net82),
    .q (net98)
  );
  dffsr_cell flop3 (
    .d (net98),
    .clk (net96),
    .s (net8),
    .r (net82),
    .q (net99)
  );
  dffsr_cell flop4 (
    .d (net99),
    .clk (net96),
    .s (net100),
    .r (net82),
    .q (net101)
  );
  dffsr_cell flop5 (
    .d (net101),
    .clk (net96),
    .s (net100),
    .r (net82),
    .q (net102)
  );
  dffsr_cell flop6 (
    .d (net102),
    .clk (net96),
    .s (net100),
    .r (net82),
    .q (net103)
  );
  dffsr_cell flop7 (
    .d (net103),
    .clk (net96),
    .s (net100),
    .r (net82),
    .q (net104)
  );
  dffsr_cell flop8 (
    .d (net104),
    .clk (net96),
    .s (net100),
    .r (net82),
    .q (net105)
  );
  dffsr_cell flop9 (
    .d (net106),
    .clk (net107),
    .s (net8),
    .r (net82),
    .q (net108)
  );
  dffsr_cell flop10 (
    .d (net108),
    .clk (net107),
    .s (net100),
    .r (net82),
    .q (net109)
  );
  dffsr_cell flop11 (
    .d (net109),
    .clk (net107),
    .s (net8),
    .r (net82),
    .q (net110)
  );
  dffsr_cell flop12 (
    .d (net110),
    .clk (net107),
    .s (net100),
    .r (net82),
    .q (net111)
  );
  dffsr_cell flop13 (
    .d (net111),
    .clk (net107),
    .s (net100),
    .r (net82),
    .q (net112)
  );
  dffsr_cell flop14 (
    .d (net112),
    .clk (net107),
    .s (net100),
    .r (net82),
    .q (net113)
  );
  dffsr_cell flop15 (
    .d (net113),
    .clk (net107),
    .s (net100),
    .r (net82),
    .q (net114)
  );
  dffsr_cell flop16 (
    .d (net114),
    .clk (net107),
    .s (net100),
    .r (net82),
    .q (net115)
  );
  mux_cell mux15 (
    .a (net116),
    .b (net117),
    .sel (net17),
    .out (net118)
  );
  mux_cell mux16 (
    .a (net119),
    .b (net117),
    .sel (net17),
    .out (net120)
  );
  mux_cell mux17 (
    .a (net117),
    .b (net116),
    .sel (net17),
    .out (net107)
  );
  mux_cell mux18 (
    .a (net117),
    .b (net119),
    .sel (net17),
    .out (net106)
  );
  mux_cell mux19 (
    .a (net121),
    .b (net117),
    .sel (net17),
    .out (net96)
  );
  mux_cell mux20 (
    .a (net122),
    .b (net117),
    .sel (net17),
    .out (net95)
  );
  mux_cell mux21 (
    .a (net117),
    .b (net121),
    .sel (net17),
    .out (net123)
  );
  mux_cell mux22 (
    .a (net117),
    .b (net122),
    .sel (net17),
    .out (net124)
  );
  mux_cell mux23 (
    .a (net125),
    .b (net117),
    .sel (net17),
    .out (net126)
  );
  mux_cell mux24 (
    .a (net127),
    .b (net117),
    .sel (net17),
    .out (net128)
  );
  mux_cell mux25 (
    .a (net117),
    .b (net125),
    .sel (net17),
    .out (net129)
  );
  mux_cell mux26 (
    .a (net117),
    .b (net127),
    .sel (net17),
    .out (net130)
  );
  mux_cell mux27 (
    .a (net131),
    .b (net117),
    .sel (net17),
    .out (net132)
  );
  mux_cell mux28 (
    .a (net133),
    .b (net117),
    .sel (net17),
    .out (net134)
  );
  mux_cell mux29 (
    .a (net117),
    .b (net131),
    .sel (net17),
    .out (net135)
  );
  mux_cell mux30 (
    .a (net117),
    .b (net133),
    .sel (net17),
    .out (net136)
  );
  mux_cell mux31 (
    .a (net137),
    .b (net117),
    .sel (net19),
    .out (net116)
  );
  mux_cell mux32 (
    .a (net138),
    .b (net117),
    .sel (net19),
    .out (net119)
  );
  mux_cell mux33 (
    .a (net117),
    .b (net137),
    .sel (net19),
    .out (net121)
  );
  mux_cell mux34 (
    .a (net117),
    .b (net138),
    .sel (net19),
    .out (net122)
  );
  mux_cell mux35 (
    .a (net139),
    .b (net117),
    .sel (net19),
    .out (net125)
  );
  mux_cell mux36 (
    .a (net140),
    .b (net117),
    .sel (net19),
    .out (net127)
  );
  mux_cell mux37 (
    .a (net117),
    .b (net139),
    .sel (net19),
    .out (net131)
  );
  mux_cell mux38 (
    .a (net117),
    .b (net140),
    .sel (net19),
    .out (net133)
  );
  mux_cell mux39 (
    .a (net4),
    .b (net117),
    .sel (net20),
    .out (net137)
  );
  mux_cell mux40 (
    .a (net5),
    .b (net117),
    .sel (net20),
    .out (net138)
  );
  mux_cell mux41 (
    .a (net117),
    .b (net4),
    .sel (net20),
    .out (net139)
  );
  mux_cell mux42 (
    .a (net117),
    .b (net5),
    .sel (net20),
    .out (net140)
  );
  dffsr_cell flop17 (
    .d (net124),
    .clk (net123),
    .s (net8),
    .r (net82),
    .q (net141)
  );
  dffsr_cell flop18 (
    .d (net141),
    .clk (net123),
    .s (net8),
    .r (net82),
    .q (net142)
  );
  dffsr_cell flop19 (
    .d (net142),
    .clk (net123),
    .s (net8),
    .r (net82),
    .q (net143)
  );
  dffsr_cell flop20 (
    .d (net143),
    .clk (net123),
    .s (net100),
    .r (net82),
    .q (net144)
  );
  dffsr_cell flop21 (
    .d (net144),
    .clk (net123),
    .s (net100),
    .r (net82),
    .q (net145)
  );
  dffsr_cell flop22 (
    .d (net145),
    .clk (net123),
    .s (net100),
    .r (net82),
    .q (net146)
  );
  dffsr_cell flop23 (
    .d (net146),
    .clk (net123),
    .s (net100),
    .r (net82),
    .q (net147)
  );
  dffsr_cell flop24 (
    .d (net147),
    .clk (net123),
    .s (net100),
    .r (net82),
    .q (net148)
  );
  dffsr_cell flop25 (
    .d (net130),
    .clk (net129),
    .s (net100),
    .r (net82),
    .q (net88)
  );
  dffsr_cell flop26 (
    .d (net88),
    .clk (net129),
    .s (net100),
    .r (net82),
    .q (net89)
  );
  dffsr_cell flop27 (
    .d (net89),
    .clk (net129),
    .s (net8),
    .r (net82),
    .q (net90)
  );
  dffsr_cell flop28 (
    .d (net90),
    .clk (net129),
    .s (net8),
    .r (net82),
    .q (net91)
  );
  dffsr_cell flop29 (
    .d (net91),
    .clk (net129),
    .s (net100),
    .r (net82),
    .q (net92)
  );
  dffsr_cell flop30 (
    .d (net92),
    .clk (net129),
    .s (net100),
    .r (net82),
    .q (net93)
  );
  dffsr_cell flop31 (
    .d (net93),
    .clk (net129),
    .s (net100),
    .r (net82),
    .q (net94)
  );
  dffsr_cell flop32 (
    .d (net94),
    .clk (net129),
    .s (net100),
    .r (net82),
    .q (net149)
  );
  dffsr_cell flop33 (
    .d (net150),
    .clk (net126),
    .s (net8),
    .r (net82),
    .q (net67)
  );
  dffsr_cell flop34 (
    .d (net67),
    .clk (net126),
    .s (net8),
    .r (net82),
    .q (net65)
  );
  dffsr_cell flop35 (
    .d (net65),
    .clk (net126),
    .s (net8),
    .r (net82),
    .q (net63)
  );
  dffsr_cell flop36 (
    .d (net63),
    .clk (net126),
    .s (net100),
    .r (net82),
    .q (net61)
  );
  dffsr_cell flop37 (
    .d (net61),
    .clk (net126),
    .s (net100),
    .r (net82),
    .q (net43)
  );
  dffsr_cell flop38 (
    .d (net43),
    .clk (net126),
    .s (net100),
    .r (net82),
    .q (net41)
  );
  dffsr_cell flop39 (
    .d (net41),
    .clk (net126),
    .s (net100),
    .r (net82),
    .q (net30)
  );
  dffsr_cell flop40 (
    .d (net128),
    .clk (net126),
    .s (net8),
    .r (net82),
    .q (net150)
  );
  dffsr_cell flop41 (
    .d (net134),
    .clk (net132),
    .s (net100),
    .r (net82),
    .q (net151)
  );
  dffsr_cell flop42 (
    .d (net151),
    .clk (net132),
    .s (net100),
    .r (net82),
    .q (net152)
  );
  dffsr_cell flop43 (
    .d (net152),
    .clk (net132),
    .s (net100),
    .r (net82),
    .q (net153)
  );
  dffsr_cell flop44 (
    .d (net153),
    .clk (net132),
    .s (net100),
    .r (net82),
    .q (net154)
  );
  dffsr_cell flop45 (
    .d (net154),
    .clk (net132),
    .s (net100),
    .r (net82),
    .q (net155)
  );
  dffsr_cell flop46 (
    .d (net155),
    .clk (net132),
    .s (net100),
    .r (net82),
    .q (net156)
  );
  dffsr_cell flop47 (
    .d (net156),
    .clk (net132),
    .s (net100),
    .r (net82),
    .q (net157)
  );
  dffsr_cell flop48 (
    .d (net157),
    .clk (net132),
    .s (net100),
    .r (net82),
    .q (net158)
  );
  dffsr_cell flop49 (
    .d (net136),
    .clk (net135),
    .s (net100),
    .r (net82),
    .q (net159)
  );
  dffsr_cell flop50 (
    .d (net159),
    .clk (net135),
    .s (net100),
    .r (net82),
    .q (net160)
  );
  dffsr_cell flop51 (
    .d (net160),
    .clk (net135),
    .s (net100),
    .r (net82),
    .q (net161)
  );
  dffsr_cell flop52 (
    .d (net161),
    .clk (net135),
    .s (net100),
    .r (net82),
    .q (net162)
  );
  dffsr_cell flop53 (
    .d (net162),
    .clk (net135),
    .s (net100),
    .r (net82),
    .q (net163)
  );
  dffsr_cell flop54 (
    .d (net163),
    .clk (net135),
    .s (net100),
    .r (net82),
    .q (net164)
  );
  dffsr_cell flop55 (
    .d (net164),
    .clk (net135),
    .s (net100),
    .r (net82),
    .q (net165)
  );
  dffsr_cell flop56 (
    .d (net165),
    .clk (net135),
    .s (net100),
    .r (net82),
    .q (net166)
  );
  dffsr_cell flop57 (
    .d (net120),
    .clk (net118),
    .s (net100),
    .r (net3),
    .q (net167)
  );
  dffsr_cell flop58 (
    .d (net167),
    .clk (net118),
    .s (net100),
    .r (net3),
    .q (net168)
  );
  dffsr_cell flop59 (
    .d (net168),
    .clk (net118),
    .s (net100),
    .r (net3),
    .q (net169)
  );
  dffsr_cell flop60 (
    .d (net169),
    .clk (net118),
    .s (net100),
    .r (net3),
    .q (net170)
  );
  dffsr_cell flop61 (
    .d (net170),
    .clk (net118),
    .s (net100),
    .r (net3),
    .q (net171)
  );
  dffsr_cell flop62 (
    .d (net171),
    .clk (net118),
    .s (net100),
    .r (net3),
    .q (net172)
  );
  dffsr_cell flop63 (
    .d (net172),
    .clk (net118),
    .s (net100),
    .r (net3),
    .q (net173)
  );
  dffsr_cell flop64 (
    .d (net173),
    .clk (net118),
    .s (net100),
    .r (net3),
    .q (net174)
  );
  dffsr_cell flop65 (
    .d (net176),
    .clk (net177),
    .s (net178),
    .r (net179),
    .q (net180),
    .notq (net176)
  );
  dffsr_cell flop66 (
    .d (net181),
    .clk (net176),
    .s (net178),
    .r (net179),
    .q (net182),
    .notq (net181)
  );
  and_cell and15 (
    .a (net183),
    .b (net184),
    .out (net185)
  );
  or_cell or2 (
    .a (net185),
    .b (net186),
    .out (net187)
  );
  or_cell or3 (
    .a (net188),
    .b (net189),
    .out (net190)
  );
  and_cell and16 (
    .a (net190),
    .b (net187),
    .out (net191)
  );
  and_cell and17 (
    .a (net180),
    .b (net192),
    .out (net186)
  );
  not_cell not2 (
    .in (net192),
    .out (net184)
  );
  not_cell not3 (
    .in (net180),
    .out (net183)
  );
  or_cell or4 (
    .a (net193),
    .b (net194),
    .out (net179)
  );
  dff_cell flop67 (
    .d (net23),
    .clk (net177),
    .q (net195)
  );
  dffsr_cell flop68 (
    .d (net196),
    .clk (net181),
    .s (net178),
    .r (net179),
    .q (net197),
    .notq (net196)
  );
  dffsr_cell flop69 (
    .d (net198),
    .clk (net196),
    .s (net178),
    .r (net179),
    .q (net199),
    .notq (net198)
  );
  dffsr_cell flop70 (
    .d (net200),
    .clk (net198),
    .s (net178),
    .r (net179),
    .q (net201),
    .notq (net200)
  );
  dffsr_cell flop71 (
    .d (net202),
    .clk (net200),
    .s (net178),
    .r (net179),
    .q (net203),
    .notq (net202)
  );
  dffsr_cell flop72 (
    .d (net204),
    .clk (net202),
    .s (net178),
    .r (net179),
    .q (net205),
    .notq (net204)
  );
  dffsr_cell flop73 (
    .d (net206),
    .clk (net204),
    .s (net178),
    .r (net179),
    .q (net207),
    .notq (net206)
  );
  mux_cell mux43 (
    .a (net98),
    .b (net99),
    .sel (net13),
    .out (net208)
  );
  mux_cell mux44 (
    .a (net97),
    .b (net98),
    .sel (net13),
    .out (net192)
  );
  and_cell and18 (
    .a (net209),
    .b (net210),
    .out (net188)
  );
  and_cell and19 (
    .a (net182),
    .b (net208),
    .out (net189)
  );
  not_cell not4 (
    .in (net208),
    .out (net210)
  );
  not_cell not5 (
    .in (net182),
    .out (net209)
  );
  and_cell and20 (
    .a (net211),
    .b (net212),
    .out (net213)
  );
  or_cell or5 (
    .a (net213),
    .b (net214),
    .out (net215)
  );
  or_cell or6 (
    .a (net216),
    .b (net217),
    .out (net218)
  );
  and_cell and21 (
    .a (net218),
    .b (net215),
    .out (net219)
  );
  and_cell and22 (
    .a (net197),
    .b (net220),
    .out (net214)
  );
  not_cell not6 (
    .in (net220),
    .out (net212)
  );
  not_cell not7 (
    .in (net197),
    .out (net211)
  );
  and_cell and23 (
    .a (net221),
    .b (net222),
    .out (net216)
  );
  and_cell and24 (
    .a (net199),
    .b (net223),
    .out (net217)
  );
  not_cell not8 (
    .in (net223),
    .out (net222)
  );
  not_cell not9 (
    .in (net199),
    .out (net221)
  );
  and_cell and25 (
    .a (net224),
    .b (net225),
    .out (net226)
  );
  or_cell or7 (
    .a (net226),
    .b (net227),
    .out (net228)
  );
  or_cell or8 (
    .a (net229),
    .b (net230),
    .out (net231)
  );
  and_cell and26 (
    .a (net231),
    .b (net228),
    .out (net232)
  );
  and_cell and27 (
    .a (net201),
    .b (net233),
    .out (net227)
  );
  not_cell not10 (
    .in (net233),
    .out (net225)
  );
  not_cell not11 (
    .in (net201),
    .out (net224)
  );
  and_cell and28 (
    .a (net234),
    .b (net235),
    .out (net229)
  );
  and_cell and29 (
    .a (net203),
    .b (net236),
    .out (net230)
  );
  not_cell not12 (
    .in (net236),
    .out (net235)
  );
  not_cell not13 (
    .in (net203),
    .out (net234)
  );
  and_cell and30 (
    .a (net237),
    .b (net238),
    .out (net239)
  );
  or_cell or9 (
    .a (net239),
    .b (net240),
    .out (net241)
  );
  or_cell or10 (
    .a (net242),
    .b (net243),
    .out (net244)
  );
  and_cell and31 (
    .a (net244),
    .b (net241),
    .out (net245)
  );
  and_cell and32 (
    .a (net205),
    .b (net246),
    .out (net240)
  );
  not_cell not14 (
    .in (net246),
    .out (net238)
  );
  not_cell not15 (
    .in (net205),
    .out (net237)
  );
  and_cell and33 (
    .a (net247),
    .b (net248),
    .out (net242)
  );
  and_cell and34 (
    .a (net207),
    .b (net249),
    .out (net243)
  );
  not_cell not16 (
    .in (net249),
    .out (net248)
  );
  not_cell not17 (
    .in (net207),
    .out (net247)
  );
  and_cell and35 (
    .a (net219),
    .b (net191),
    .out (net250)
  );
  and_cell and36 (
    .a (net232),
    .b (net250),
    .out (net251)
  );
  and_cell and37 (
    .a (net245),
    .b (net251),
    .out (net23)
  );
  mux_cell mux45 (
    .a (net101),
    .b (net102),
    .sel (net13),
    .out (net223)
  );
  mux_cell mux46 (
    .a (net99),
    .b (net101),
    .sel (net13),
    .out (net220)
  );
  mux_cell mux47 (
    .a (net103),
    .b (net104),
    .sel (net13),
    .out (net236)
  );
  mux_cell mux48 (
    .a (net102),
    .b (net103),
    .sel (net13),
    .out (net233)
  );
  mux_cell mux49 (
    .a (net105),
    .b (net252),
    .sel (net13),
    .out (net249)
  );
  mux_cell mux50 (
    .a (net104),
    .b (net105),
    .sel (net13),
    .out (net246)
  );
  dffsr_cell flop74 (
    .d (net13),
    .clk (net195),
    .s (net178),
    .r (net179),
    .q (net253),
    .notq (net13)
  );
  and_cell and38 (
    .a (net253),
    .b (net23),
    .out (net254)
  );
  dff_cell flop75 (
    .d (net254),
    .clk (net177),
    .q (net194)
  );
  dffsr_cell flop76 (
    .d (net255),
    .clk (net13),
    .s (net256),
    .r (net257),
    .q (net258),
    .notq (net255)
  );
  dffsr_cell flop77 (
    .d (net259),
    .clk (net255),
    .s (net256),
    .r (net257),
    .q (net260),
    .notq (net259)
  );
  and_cell and39 (
    .a (net261),
    .b (net262),
    .out (net263)
  );
  or_cell or11 (
    .a (net263),
    .b (net264),
    .out (net265)
  );
  or_cell or12 (
    .a (net266),
    .b (net267),
    .out (net268)
  );
  and_cell and40 (
    .a (net268),
    .b (net265),
    .out (net269)
  );
  and_cell and41 (
    .a (net258),
    .b (net270),
    .out (net264)
  );
  not_cell not18 (
    .in (net270),
    .out (net262)
  );
  not_cell not19 (
    .in (net258),
    .out (net261)
  );
  or_cell or13 (
    .a (net193),
    .b (net271),
    .out (net257)
  );
  dff_cell flop78 (
    .d (net22),
    .clk (net13),
    .q (net272)
  );
  dffsr_cell flop79 (
    .d (net273),
    .clk (net259),
    .s (net256),
    .r (net257),
    .q (net274),
    .notq (net273)
  );
  dffsr_cell flop80 (
    .d (net275),
    .clk (net273),
    .s (net256),
    .r (net257),
    .q (net276),
    .notq (net275)
  );
  dffsr_cell flop81 (
    .d (net277),
    .clk (net275),
    .s (net256),
    .r (net257),
    .q (net278),
    .notq (net277)
  );
  dffsr_cell flop82 (
    .d (net279),
    .clk (net277),
    .s (net256),
    .r (net257),
    .q (net280),
    .notq (net279)
  );
  dffsr_cell flop83 (
    .d (net281),
    .clk (net279),
    .s (net256),
    .r (net257),
    .q (net282),
    .notq (net281)
  );
  dffsr_cell flop84 (
    .d (net283),
    .clk (net281),
    .s (net256),
    .r (net257),
    .q (net284),
    .notq (net283)
  );
  mux_cell mux51 (
    .a (net142),
    .b (net143),
    .sel (net285),
    .out (net286)
  );
  mux_cell mux52 (
    .a (net141),
    .b (net142),
    .sel (net285),
    .out (net270)
  );
  and_cell and42 (
    .a (net287),
    .b (net288),
    .out (net266)
  );
  and_cell and43 (
    .a (net260),
    .b (net286),
    .out (net267)
  );
  not_cell not20 (
    .in (net286),
    .out (net288)
  );
  not_cell not21 (
    .in (net260),
    .out (net287)
  );
  and_cell and44 (
    .a (net289),
    .b (net290),
    .out (net291)
  );
  or_cell or14 (
    .a (net291),
    .b (net292),
    .out (net293)
  );
  or_cell or15 (
    .a (net294),
    .b (net295),
    .out (net296)
  );
  and_cell and45 (
    .a (net296),
    .b (net293),
    .out (net297)
  );
  and_cell and46 (
    .a (net274),
    .b (net298),
    .out (net292)
  );
  not_cell not22 (
    .in (net298),
    .out (net290)
  );
  not_cell not23 (
    .in (net274),
    .out (net289)
  );
  and_cell and47 (
    .a (net299),
    .b (net300),
    .out (net294)
  );
  and_cell and48 (
    .a (net276),
    .b (net301),
    .out (net295)
  );
  not_cell not24 (
    .in (net301),
    .out (net300)
  );
  not_cell not25 (
    .in (net276),
    .out (net299)
  );
  and_cell and49 (
    .a (net302),
    .b (net303),
    .out (net304)
  );
  or_cell or16 (
    .a (net304),
    .b (net305),
    .out (net306)
  );
  or_cell or17 (
    .a (net307),
    .b (net308),
    .out (net309)
  );
  and_cell and50 (
    .a (net309),
    .b (net306),
    .out (net310)
  );
  and_cell and51 (
    .a (net278),
    .b (net311),
    .out (net305)
  );
  not_cell not26 (
    .in (net311),
    .out (net303)
  );
  not_cell not27 (
    .in (net278),
    .out (net302)
  );
  and_cell and52 (
    .a (net312),
    .b (net313),
    .out (net307)
  );
  and_cell and53 (
    .a (net280),
    .b (net314),
    .out (net308)
  );
  not_cell not28 (
    .in (net314),
    .out (net313)
  );
  not_cell not29 (
    .in (net280),
    .out (net312)
  );
  and_cell and54 (
    .a (net315),
    .b (net316),
    .out (net317)
  );
  or_cell or18 (
    .a (net317),
    .b (net318),
    .out (net319)
  );
  or_cell or19 (
    .a (net320),
    .b (net321),
    .out (net322)
  );
  and_cell and55 (
    .a (net322),
    .b (net319),
    .out (net323)
  );
  and_cell and56 (
    .a (net282),
    .b (net324),
    .out (net318)
  );
  not_cell not30 (
    .in (net324),
    .out (net316)
  );
  not_cell not31 (
    .in (net282),
    .out (net315)
  );
  and_cell and57 (
    .a (net325),
    .b (net326),
    .out (net320)
  );
  and_cell and58 (
    .a (net284),
    .b (net327),
    .out (net321)
  );
  not_cell not32 (
    .in (net327),
    .out (net326)
  );
  not_cell not33 (
    .in (net284),
    .out (net325)
  );
  and_cell and59 (
    .a (net297),
    .b (net269),
    .out (net328)
  );
  and_cell and60 (
    .a (net310),
    .b (net328),
    .out (net329)
  );
  and_cell and61 (
    .a (net323),
    .b (net329),
    .out (net22)
  );
  mux_cell mux53 (
    .a (net144),
    .b (net145),
    .sel (net285),
    .out (net301)
  );
  mux_cell mux54 (
    .a (net143),
    .b (net144),
    .sel (net285),
    .out (net298)
  );
  mux_cell mux55 (
    .a (net146),
    .b (net147),
    .sel (net285),
    .out (net314)
  );
  mux_cell mux56 (
    .a (net145),
    .b (net146),
    .sel (net285),
    .out (net311)
  );
  mux_cell mux57 (
    .a (net148),
    .b (net330),
    .sel (net285),
    .out (net327)
  );
  mux_cell mux58 (
    .a (net147),
    .b (net148),
    .sel (net285),
    .out (net324)
  );
  dffsr_cell flop85 (
    .d (net285),
    .clk (net272),
    .s (net256),
    .r (net257),
    .q (net331),
    .notq (net285)
  );
  and_cell and62 (
    .a (net331),
    .b (net22),
    .out (net332)
  );
  dff_cell flop86 (
    .d (net332),
    .clk (net13),
    .q (net271),
    .notq (net14)
  );
  dffsr_cell flop87 (
    .d (net167),
    .clk (net334),
    .s (net333),
    .r (net3),
    .q (net17)
  );
  dffsr_cell flop88 (
    .d (net168),
    .clk (net334),
    .s (net333),
    .r (net3),
    .q (net19)
  );
  dffsr_cell flop89 (
    .d (net169),
    .clk (net334),
    .s (net333),
    .r (net3),
    .q (net20)
  );
  not_cell not34 (
    .in (net4),
    .out (net335)
  );
  dffsr_cell flop90 (
    .d (net174),
    .clk (net335),
    .r (net3),
    .q (net334)
  );
  not_cell not35 (
    .in (net6),
    .out (net193)
  );
  dffsr_cell flop91 (
    .d (net28),
    .clk (net16),
    .s (net193),
    .r (net336),
    .q (net29),
    .notq (net80)
  );
  dffsr_cell flop92 (
    .d (net27),
    .clk (net16),
    .s (net193),
    .r (net336),
    .q (net40),
    .notq (net78)
  );
  dffsr_cell flop93 (
    .d (net35),
    .clk (net16),
    .s (net193),
    .r (net336),
    .q (net42),
    .notq (net76)
  );
  dffsr_cell flop94 (
    .d (net39),
    .clk (net16),
    .s (net193),
    .r (net336),
    .q (net60),
    .notq (net74)
  );
  dffsr_cell flop95 (
    .d (net47),
    .clk (net16),
    .s (net193),
    .r (net336),
    .q (net62),
    .notq (net72)
  );
  dffsr_cell flop96 (
    .d (net51),
    .clk (net16),
    .s (net193),
    .r (net336),
    .q (net64),
    .notq (net70)
  );
  dffsr_cell flop97 (
    .d (net55),
    .clk (net16),
    .s (net193),
    .r (net336),
    .q (net66),
    .notq (net68)
  );
  dffsr_cell flop98 (
    .d (net59),
    .clk (net16),
    .s (net193),
    .r (net336),
    .q (net31),
    .notq (net337)
  );
  or_cell or20 (
    .a (net1),
    .b (net21),
    .out (net15)
  );
  dffsr_cell flop99 (
    .d (net338),
    .clk (net339),
    .s (net340),
    .r (net193),
    .q (net21)
  );
  not_cell not36 (
    .in (net331),
    .out (net339)
  );
  xor_cell xor8 (
    .a (net343),
    .b (net31),
    .out (net10)
  );
  xor_cell xor9 (
    .a (net337),
    .b (net343),
    .out (net11)
  );
  xor_cell xor10 (
    .a (net66),
    .b (net343),
    .out (net9)
  );
  xor_cell xor11 (
    .a (net343),
    .b (net68),
    .out (net12)
  );
  dff_cell flop100 (
    .d (net7),
    .clk (net13),
    .q (net343)
  );
  mux_cell mux59 (
    .a (net344),
    .b (net345),
    .sel (net109),
    .out (net346)
  );
  dff_cell flop101 (
    .d (net347),
    .clk (net15),
    .q (net348),
    .notq (net347)
  );
  dff_cell flop102 (
    .d (net349),
    .clk (net344),
    .q (net350),
    .notq (net349)
  );
  mux_cell mux60 (
    .a (net346),
    .b (net351),
    .sel (net110),
    .out (net16)
  );
  mux_cell mux61 (
    .a (net15),
    .b (net348),
    .sel (net108),
    .out (net344)
  );
  dff_cell flop103 (
    .d (net352),
    .clk (net350),
    .q (net345),
    .notq (net352)
  );
  dff_cell flop104 (
    .d (net353),
    .clk (net346),
    .q (net354),
    .notq (net353)
  );
  dff_cell flop105 (
    .d (net355),
    .clk (net354),
    .q (net356),
    .notq (net355)
  );
  dff_cell flop106 (
    .d (net357),
    .clk (net356),
    .q (net358),
    .notq (net357)
  );
  dff_cell flop107 (
    .d (net359),
    .clk (net358),
    .q (net351),
    .notq (net359)
  );
  and_cell and63 (
    .a (net64),
    .b (net360),
    .out (net361)
  );
  and_cell and64 (
    .a (net66),
    .b (net31),
    .out (net360)
  );
  and_cell and65 (
    .a (net60),
    .b (net362),
    .out (net363)
  );
  and_cell and66 (
    .a (net62),
    .b (net361),
    .out (net362)
  );
  and_cell and67 (
    .a (net35),
    .b (net363),
    .out (net364)
  );
  and_cell and68 (
    .a (net29),
    .b (net365),
    .out (net366)
  );
  and_cell and69 (
    .a (net40),
    .b (net364),
    .out (net365)
  );
  dff_cell flop108 (
    .d (net366),
    .clk (net16),
    .q (net177)
  );
endmodule
