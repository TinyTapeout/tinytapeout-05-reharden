/* Automatically generated from https://wokwi.com/projects/380361576213660673 */

`default_nettype none

module tt_um_wokwi_380361576213660673(
  input  wire [7:0] ui_in,    // Dedicated inputs
  output wire [7:0] uo_out,    // Dedicated outputs
  input  wire [7:0] uio_in,    // IOs: Input path
  output wire [7:0] uio_out,    // IOs: Output path
  output wire [7:0] uio_oe,    // IOs: Enable path (active high: 0=input, 1=output)
  input ena,
  input clk,
  input rst_n
);
  wire net1 = clk;
  wire net2 = rst_n;
  wire net3 = ui_in[0];
  wire net4 = ui_in[1];
  wire net5 = ui_in[2];
  wire net6 = ui_in[3];
  wire net7 = ui_in[4];
  wire net8 = ui_in[5];
  wire net9 = ui_in[6];
  wire net10 = ui_in[7];
  wire net11;
  wire net12;
  wire net13;
  wire net14;
  wire net15;
  wire net16;
  wire net17;
  wire net18;
  wire net19 = uio_in[0];
  wire net20 = 1'b0;
  wire net21 = uio_in[1];
  wire net22 = 1'b0;
  wire net23 = 1'b1;
  wire net24 = uio_in[4];
  wire net25 = 1'b0;
  wire net26 = uio_in[5];
  wire net27 = 1'b0;
  wire net28 = uio_in[6];
  wire net29 = 1'b0;
  wire net30 = uio_in[7];
  wire net31 = 1'b0;
  wire net32;
  wire net33;
  wire net34;
  wire net35;
  wire net36;
  wire net37;
  wire net38;
  wire net39;
  wire net40;
  wire net41;
  wire net42;
  wire net43;
  wire net44;
  wire net45;
  wire net46;
  wire net47;
  wire net48;
  wire net49;
  wire net50;
  wire net51;
  wire net52;
  wire net53;
  wire net54;
  wire net55;
  wire net56;
  wire net57;
  wire net58;
  wire net59;
  wire net60;
  wire net61;
  wire net62;
  wire net63;
  wire net64;
  wire net65;
  wire net66;
  wire net67;
  wire net68;
  wire net69;
  wire net70;
  wire net71;
  wire net72;
  wire net73;
  wire net74;
  wire net75;
  wire net76;
  wire net77;
  wire net78;
  wire net79;
  wire net80;
  wire net81;
  wire net82;
  wire net83;
  wire net84;
  wire net85;
  wire net86;
  wire net87;
  wire net88;
  wire net89;
  wire net90;
  wire net91;
  wire net92;
  wire net93;
  wire net94;
  wire net95;
  wire net96;
  wire net97;
  wire net98;
  wire net99;
  wire net100;
  wire net101;
  wire net102;
  wire net103 = 1'b0;
  wire net104;
  wire net105;
  wire net106;
  wire net107;
  wire net108;
  wire net109;
  wire net110;
  wire net111 = 1'b0;
  wire net112;
  wire net113;
  wire net114;
  wire net115;
  wire net116;
  wire net117;
  wire net118 = 1'b0;
  wire net119;
  wire net120;
  wire net121;
  wire net122;
  wire net123;
  wire net124;
  wire net125;
  wire net126;
  wire net127;
  wire net128;
  wire net129;
  wire net130;
  wire net131;
  wire net132;
  wire net133;
  wire net134;
  wire net135;
  wire net136;
  wire net137;
  wire net138;
  wire net139;
  wire net140;
  wire net141;
  wire net142;
  wire net143;
  wire net144;
  wire net145;
  wire net146;
  wire net147;
  wire net148;
  wire net149;
  wire net150;
  wire net151;
  wire net152;
  wire net153;
  wire net154;
  wire net155;
  wire net156;
  wire net157;
  wire net158;
  wire net159;
  wire net160;
  wire net161;
  wire net162;
  wire net163;
  wire net164;
  wire net165;
  wire net166;
  wire net167;
  wire net168 = 1'b0;
  wire net169;
  wire net170;
  wire net171;
  wire net172;
  wire net173;
  wire net174;
  wire net175;
  wire net176;
  wire net177;
  wire net178;
  wire net179;
  wire net180;
  wire net181;
  wire net182;
  wire net183;
  wire net184;
  wire net185;
  wire net186;
  wire net187;
  wire net188;
  wire net189;
  wire net190;
  wire net191;
  wire net192;
  wire net193;
  wire net194;
  wire net195;
  wire net196;
  wire net197;
  wire net198;
  wire net199;
  wire net200;
  wire net201;
  wire net202;
  wire net203;
  wire net204;
  wire net205 = 1'b0;
  wire net206;
  wire net207;
  wire net208;
  wire net209;
  wire net210;
  wire net211;
  wire net212;
  wire net213;
  wire net214;
  wire net215;
  wire net216;
  wire net217;
  wire net218;
  wire net219;
  wire net220;
  wire net221;
  wire net222;
  wire net223;
  wire net224;
  wire net225;
  wire net226;
  wire net227;
  wire net228;
  wire net229;
  wire net230;
  wire net231;
  wire net232;
  wire net233;
  wire net234;
  wire net235;
  wire net236 = 1'b0;
  wire net237;
  wire net238;
  wire net239;
  wire net240;
  wire net241;
  wire net242;
  wire net243;
  wire net244;
  wire net245;
  wire net246;
  wire net247;
  wire net248;
  wire net249;
  wire net250;
  wire net251;
  wire net252;
  wire net253;
  wire net254;
  wire net255;
  wire net256;
  wire net257;
  wire net258;
  wire net259;
  wire net260;
  wire net261;
  wire net262;
  wire net263;
  wire net264;
  wire net265;
  wire net266;
  wire net267;
  wire net268;
  wire net269;
  wire net270;
  wire net271;
  wire net272;
  wire net273;
  wire net274;
  wire net275;
  wire net276;
  wire net277;
  wire net278;
  wire net279;
  wire net280;
  wire net281;
  wire net282;
  wire net283;
  wire net284;
  wire net285;
  wire net286 = 1'b1;
  wire net287;
  wire net288;
  wire net289 = 1'b0;
  wire net290;
  wire net291;
  wire net292;
  wire net293;
  wire net294 = 1'b0;
  wire net295;
  wire net296;
  wire net297;
  wire net298;
  wire net299;
  wire net300;
  wire net301;
  wire net302;
  wire net303;
  wire net304;
  wire net305;
  wire net306;
  wire net307;
  wire net308;
  wire net309;
  wire net310;
  wire net311;
  wire net312;
  wire net313;
  wire net314;
  wire net315;
  wire net316;
  wire net317;
  wire net318;
  wire net319;
  wire net320;
  wire net321;
  wire net322;
  wire net323;
  wire net324;
  wire net325;
  wire net326;
  wire net327;
  wire net328;
  wire net329;
  wire net330;
  wire net331;
  wire net332;
  wire net333;
  wire net334;
  wire net335;
  wire net336;
  wire net337;
  wire net338;
  wire net339 = 1'b0;
  wire net340;
  wire net341;
  wire net342;
  wire net343;
  wire net344;
  wire net345;
  wire net346;
  wire net347;
  wire net348;
  wire net349;
  wire net350;
  wire net351;
  wire net352;
  wire net353;
  wire net354;
  wire net355;
  wire net356;
  wire net357;
  wire net358;
  wire net359;
  wire net360;
  wire net361 = 1'b0;
  wire net362;
  wire net363;
  wire net364;
  wire net365;
  wire net366;
  wire net367;
  wire net368;
  wire net369;
  wire net370;
  wire net371;
  wire net372;
  wire net373;
  wire net374;
  wire net375;
  wire net376;
  wire net377;
  wire net378;
  wire net379;
  wire net380;
  wire net381;
  wire net382;
  wire net383;
  wire net384;
  wire net385;
  wire net386;
  wire net387;
  wire net388;
  wire net389;
  wire net390;
  wire net391;
  wire net392;
  wire net393;
  wire net394;
  wire net395;
  wire net396 = 1'b0;
  wire net397;
  wire net398;
  wire net399;
  wire net400;
  wire net401;
  wire net402;
  wire net403;
  wire net404;
  wire net405;
  wire net406;
  wire net407;
  wire net408;
  wire net409;
  wire net410;
  wire net411;
  wire net412;
  wire net413;
  wire net414;
  wire net415;
  wire net416;
  wire net417;
  wire net418;
  wire net419;
  wire net420;
  wire net421;
  wire net422 = 1'b1;
  wire net423;
  wire net424;
  wire net425;
  wire net426;
  wire net427;
  wire net428;
  wire net429;
  wire net430;
  wire net431;
  wire net432;
  wire net433 = 1'b0;
  wire net434;
  wire net435;
  wire net436;
  wire net437;
  wire net438;
  wire net439;
  wire net440;
  wire net441;
  wire net442;
  wire net443;
  wire net444;
  wire net445;
  wire net446;
  wire net447;
  wire net448;
  wire net449;
  wire net450;
  wire net451;
  wire net452;
  wire net453;
  wire net454;
  wire net455;
  wire net456 = 1'b1;
  wire net457 = 1'b0;
  wire net458;
  wire net459;
  wire net460;
  wire net461;
  wire net462;
  wire net463;
  wire net464;
  wire net465;
  wire net466;
  wire net467;
  wire net468;
  wire net469;
  wire net470;
  wire net471;
  wire net472;
  wire net473;
  wire net474;
  wire net475;
  wire net476;
  wire net477;
  wire net478;
  wire net479;
  wire net480;
  wire net481;
  wire net482;
  wire net483;
  wire net484;
  wire net485;
  wire net486;
  wire net487;
  wire net488;
  wire net489;
  wire net490 = 1'b1;
  wire net491;
  wire net492;
  wire net493;
  wire net494;
  wire net495;
  wire net496 = 1'b0;
  wire net497;
  wire net498;
  wire net499;
  wire net500;
  wire net501;
  wire net502;
  wire net503;
  wire net504;
  wire net505;
  wire net506;
  wire net507;
  wire net508;
  wire net509;
  wire net510;
  wire net511;
  wire net512;
  wire net513;
  wire net514;
  wire net515;
  wire net516;
  wire net517;
  wire net518;
  wire net519;
  wire net520;
  wire net521;
  wire net522;
  wire net523;
  wire net524;
  wire net525;
  wire net526 = 1'b1;
  wire net527 = 1'b0;
  wire net528;
  wire net529;
  wire net530;
  wire net531;
  wire net532;
  wire net533;
  wire net534;
  wire net535;
  wire net536;
  wire net537;
  wire net538;
  wire net539;
  wire net540;
  wire net541;
  wire net542;
  wire net543;
  wire net544;
  wire net545;
  wire net546;
  wire net547;
  wire net548;
  wire net549;
  wire net550;
  wire net551;
  wire net552;
  wire net553;
  wire net554;
  wire net555;
  wire net556;
  wire net557;
  wire net558;
  wire net559;
  wire net560 = 1'b1;
  wire net561;
  wire net562;
  wire net563;
  wire net564;
  wire net565;
  wire net566 = 1'b0;
  wire net567;
  wire net568;
  wire net569;
  wire net570;
  wire net571;
  wire net572;
  wire net573;
  wire net574;
  wire net575;
  wire net576;
  wire net577;
  wire net578;
  wire net579;
  wire net580;
  wire net581;
  wire net582;
  wire net583;
  wire net584;
  wire net585;
  wire net586;
  wire net587;
  wire net588;
  wire net589;
  wire net590;
  wire net591;
  wire net592;
  wire net593;
  wire net594;
  wire net595;
  wire net596 = 1'b1;
  wire net597;
  wire net598;
  wire net599;
  wire net600;
  wire net601;
  wire net602;
  wire net603;
  wire net604;
  wire net605;
  wire net606;
  wire net607 = 1'b0;
  wire net608;
  wire net609;
  wire net610;
  wire net611;
  wire net612;
  wire net613;
  wire net614;
  wire net615;
  wire net616;
  wire net617;
  wire net618;
  wire net619;
  wire net620;
  wire net621;
  wire net622;
  wire net623;
  wire net624;
  wire net625;
  wire net626;
  wire net627;
  wire net628;
  wire net629;
  wire net630;
  wire net631;
  wire net632;
  wire net633;
  wire net634;
  wire net635;
  wire net636;
  wire net637;
  wire net638;
  wire net639 = 1'b0;
  wire net640;
  wire net641;
  wire net642;
  wire net643;
  wire net644;
  wire net645;
  wire net646;
  wire net647;
  wire net648;
  wire net649;
  wire net650;
  wire net651;
  wire net652;
  wire net653;
  wire net654;
  wire net655;
  wire net656;
  wire net657;
  wire net658;
  wire net659;
  wire net660;
  wire net661;
  wire net662;
  wire net663;
  wire net664;
  wire net665;
  wire net666;
  wire net667;
  wire net668;
  wire net669;
  wire net670;
  wire net671;
  wire net672;
  wire net673;
  wire net674;
  wire net675;
  wire net676;
  wire net677;
  wire net678;
  wire net679;
  wire net680;
  wire net681;
  wire net682;
  wire net683;
  wire net684;
  wire net685;
  wire net686;
  wire net687;
  wire net688;
  wire net689;
  wire net690;
  wire net691;
  wire net692;
  wire net693;
  wire net694;
  wire net695;
  wire net696;
  wire net697;
  wire net698;
  wire net699;
  wire net700;
  wire net701;
  wire net702;
  wire net703;
  wire net704;
  wire net705;
  wire net706;
  wire net707;
  wire net708;
  wire net709;
  wire net710;
  wire net711;
  wire net712;
  wire net713;
  wire net714;
  wire net715;
  wire net716;
  wire net717;
  wire net718;
  wire net719;
  wire net720;
  wire net721;
  wire net722;
  wire net723;
  wire net724;
  wire net725;
  wire net726;
  wire net727;
  wire net728;
  wire net729;
  wire net730;
  wire net731;
  wire net732;
  wire net733;
  wire net734;
  wire net735;
  wire net736;
  wire net737;
  wire net738;
  wire net739;
  wire net740;
  wire net741;
  wire net742;
  wire net743;
  wire net744;
  wire net745;
  wire net746;
  wire net747;
  wire net748;
  wire net749;
  wire net750;
  wire net751;
  wire net752;
  wire net753;
  wire net754;
  wire net755;
  wire net756;
  wire net757;
  wire net758;
  wire net759;
  wire net760;
  wire net761;
  wire net762;
  wire net763;
  wire net764;
  wire net765;
  wire net766;
  wire net767;
  wire net768;
  wire net769;
  wire net770;
  wire net771;
  wire net772;
  wire net773;
  wire net774;
  wire net775;
  wire net776;
  wire net777;
  wire net778;
  wire net779;
  wire net780;
  wire net781;
  wire net782;
  wire net783;
  wire net784;
  wire net785;
  wire net786;
  wire net787;
  wire net788;
  wire net789;
  wire net790;
  wire net791;
  wire net792;
  wire net793;
  wire net794;
  wire net795;
  wire net796;
  wire net797;
  wire net798;
  wire net799;
  wire net800;
  wire net801;
  wire net802;
  wire net803;
  wire net804;
  wire net805;
  wire net806;
  wire net807;
  wire net808;
  wire net809;
  wire net810;
  wire net811;
  wire net812;
  wire net813;

  assign uo_out[0] = net11;
  assign uo_out[1] = net12;
  assign uo_out[2] = net13;
  assign uo_out[3] = net14;
  assign uo_out[4] = net15;
  assign uo_out[5] = net16;
  assign uo_out[6] = net17;
  assign uo_out[7] = net18;
  assign uio_out[0] = net20;
  assign uio_oe[0] = net20;
  assign uio_out[1] = net20;
  assign uio_oe[1] = net20;
  assign uio_out[2] = net22;
  assign uio_oe[2] = net23;
  assign uio_out[3] = net22;
  assign uio_oe[3] = net23;
  assign uio_out[4] = 0;
  assign uio_oe[4] = net25;
  assign uio_out[5] = net27;
  assign uio_oe[5] = net27;
  assign uio_out[6] = net29;
  assign uio_oe[6] = net29;
  assign uio_out[7] = net31;
  assign uio_oe[7] = net31;

  not_cell not1 (
    .in (net32),
    .out (net33)
  );
  not_cell not2 (
    .in (net34),
    .out (net35)
  );
  dff_cell flop5 (
    .d (net36),
    .clk (net24),
    .q (net34),
    .notq (net37)
  );
  dff_cell flop6 (
    .d (net38),
    .clk (net24),
    .q (net32),
    .notq (net39)
  );
  and_cell and55 (
    .a (net32),
    .b (net37),
    .out (net36)
  );
  and_cell and56 (
    .a (net39),
    .b (net37),
    .out (net38)
  );
  and_cell and1 (
    .a (net32),
    .b (net35),
    .out (net40)
  );
  and_cell and3 (
    .a (net33),
    .b (net35),
    .out (net41)
  );
  and_cell and2 (
    .a (net41),
    .b (net42),
    .out (net43)
  );
  and_cell and4 (
    .a (net40),
    .b (net44),
    .out (net45)
  );
  and_cell and5 (
    .a (net46),
    .b (net47),
    .out (net48)
  );
  or_cell or1 (
    .a (net43),
    .b (net45),
    .out (net49)
  );
  or_cell or2 (
    .a (net49),
    .b (net48),
    .out (net50)
  );
  and_cell and6 (
    .a (net41),
    .b (net51),
    .out (net52)
  );
  and_cell and7 (
    .a (net40),
    .b (net53),
    .out (net54)
  );
  and_cell and8 (
    .a (net46),
    .b (net55),
    .out (net56)
  );
  or_cell or3 (
    .a (net52),
    .b (net54),
    .out (net57)
  );
  or_cell or4 (
    .a (net57),
    .b (net56),
    .out (net58)
  );
  and_cell and9 (
    .a (net41),
    .b (net59),
    .out (net60)
  );
  and_cell and10 (
    .a (net40),
    .b (net61),
    .out (net62)
  );
  and_cell and11 (
    .a (net46),
    .b (net63),
    .out (net64)
  );
  or_cell or5 (
    .a (net60),
    .b (net62),
    .out (net65)
  );
  or_cell or6 (
    .a (net65),
    .b (net64),
    .out (net66)
  );
  and_cell and12 (
    .a (net41),
    .b (net67),
    .out (net68)
  );
  and_cell and13 (
    .a (net40),
    .b (net69),
    .out (net70)
  );
  and_cell and14 (
    .a (net46),
    .b (net71),
    .out (net72)
  );
  or_cell or7 (
    .a (net68),
    .b (net70),
    .out (net73)
  );
  or_cell or8 (
    .a (net73),
    .b (net72),
    .out (net74)
  );
  and_cell and15 (
    .a (net41),
    .b (net75),
    .out (net76)
  );
  and_cell and16 (
    .a (net40),
    .b (net77),
    .out (net78)
  );
  and_cell and17 (
    .a (net46),
    .b (net79),
    .out (net80)
  );
  or_cell or9 (
    .a (net76),
    .b (net78),
    .out (net81)
  );
  or_cell or10 (
    .a (net81),
    .b (net80),
    .out (net11)
  );
  and_cell and18 (
    .a (net41),
    .b (net82),
    .out (net83)
  );
  and_cell and19 (
    .a (net40),
    .b (net84),
    .out (net85)
  );
  and_cell and20 (
    .a (net46),
    .b (net86),
    .out (net87)
  );
  or_cell or11 (
    .a (net83),
    .b (net85),
    .out (net88)
  );
  or_cell or12 (
    .a (net88),
    .b (net87),
    .out (net12)
  );
  and_cell and21 (
    .a (net41),
    .b (net89),
    .out (net90)
  );
  and_cell and22 (
    .a (net40),
    .b (net91),
    .out (net92)
  );
  and_cell and23 (
    .a (net46),
    .b (net93),
    .out (net94)
  );
  or_cell or13 (
    .a (net90),
    .b (net92),
    .out (net95)
  );
  or_cell or14 (
    .a (net95),
    .b (net94),
    .out (net13)
  );
  and_cell and24 (
    .a (net41),
    .b (net96),
    .out (net97)
  );
  and_cell and25 (
    .a (net40),
    .b (net98),
    .out (net99)
  );
  and_cell and26 (
    .a (net46),
    .b (net100),
    .out (net101)
  );
  or_cell or15 (
    .a (net97),
    .b (net99),
    .out (net102)
  );
  or_cell or16 (
    .a (net102),
    .b (net101),
    .out (net14)
  );
  and_cell and27 (
    .a (net41),
    .b (net103),
    .out (net104)
  );
  and_cell and28 (
    .a (net40),
    .b (net105),
    .out (net106)
  );
  and_cell and29 (
    .a (net46),
    .b (net107),
    .out (net108)
  );
  or_cell or17 (
    .a (net104),
    .b (net106),
    .out (net109)
  );
  or_cell or18 (
    .a (net109),
    .b (net108),
    .out (net15)
  );
  and_cell and30 (
    .a (net33),
    .b (net34),
    .out (net46)
  );
  dffsr_cell flop18 (
    .d (net110),
    .clk (net1),
    .s (net111),
    .r (net112),
    .q (net113)
  );
  dffsr_cell flop19 (
    .d (net114),
    .clk (net1),
    .s (net111),
    .r (net112),
    .q (net115)
  );
  dffsr_cell flop11 (
    .d (net116),
    .clk (net1),
    .s (net117),
    .r (net118),
    .q (net42),
    .notq (net119)
  );
  mux_cell mux1 (
    .a (net42),
    .b (net119),
    .sel (net120),
    .out (net121)
  );
  xor_cell xor1 (
    .a (net51),
    .b (net121),
    .out (net122)
  );
  dffsr_cell flop12 (
    .d (net123),
    .clk (net1),
    .s (net118),
    .r (net117),
    .q (net51),
    .notq (net124)
  );
  and_cell and67 (
    .a (net42),
    .b (net51),
    .out (net125)
  );
  and_cell and68 (
    .a (net124),
    .b (net119),
    .out (net126)
  );
  mux_cell mux2 (
    .a (net125),
    .b (net126),
    .sel (net120),
    .out (net127)
  );
  xor_cell xor2 (
    .a (net59),
    .b (net127),
    .out (net128)
  );
  dffsr_cell flop13 (
    .d (net129),
    .clk (net1),
    .s (net118),
    .r (net117),
    .q (net59),
    .notq (net130)
  );
  and_cell and69 (
    .a (net125),
    .b (net59),
    .out (net131)
  );
  and_cell and70 (
    .a (net130),
    .b (net126),
    .out (net132)
  );
  mux_cell mux3 (
    .a (net131),
    .b (net132),
    .sel (net120),
    .out (net133)
  );
  xor_cell xor3 (
    .a (net67),
    .b (net133),
    .out (net134)
  );
  dffsr_cell flop14 (
    .d (net135),
    .clk (net1),
    .s (net117),
    .r (net118),
    .q (net67),
    .notq (net136)
  );
  not_cell not15 (
    .in (net137),
    .out (net117)
  );
  and_cell and71 (
    .a (net138),
    .b (net139),
    .out (net140)
  );
  and_cell and72 (
    .a (net59),
    .b (net67),
    .out (net141)
  );
  and_cell and73 (
    .a (net51),
    .b (net141),
    .out (net142)
  );
  and_cell and74 (
    .a (net143),
    .b (net142),
    .out (net144)
  );
  nand_cell nand7 (
    .a (net42),
    .b (net144),
    .out (net138)
  );
  not_cell not16 (
    .in (net120),
    .out (net143)
  );
  nand_cell nand8 (
    .a (net119),
    .b (net145),
    .out (net139)
  );
  and_cell and75 (
    .a (net120),
    .b (net146),
    .out (net145)
  );
  and_cell and76 (
    .a (net124),
    .b (net147),
    .out (net146)
  );
  and_cell and77 (
    .a (net59),
    .b (net136),
    .out (net147)
  );
  and_cell and78 (
    .a (net140),
    .b (net148),
    .out (net149)
  );
  or_cell or27 (
    .a (net113),
    .b (net115),
    .out (net150)
  );
  nand_cell nand9 (
    .a (net113),
    .b (net115),
    .out (net151)
  );
  and_cell and79 (
    .a (net150),
    .b (net151),
    .out (net152)
  );
  and_cell and80 (
    .a (net152),
    .b (net26),
    .out (net148)
  );
  and_cell and81 (
    .a (net153),
    .b (net115),
    .out (net120)
  );
  not_cell not17 (
    .in (net113),
    .out (net153)
  );
  dffsr_cell flop1 (
    .d (net154),
    .clk (net1),
    .s (net111),
    .r (net112),
    .q (net155)
  );
  dffsr_cell flop2 (
    .d (net156),
    .clk (net1),
    .s (net111),
    .r (net112),
    .q (net157)
  );
  dffsr_cell flop3 (
    .d (net158),
    .clk (net1),
    .s (net111),
    .r (net112),
    .q (net159)
  );
  dffsr_cell flop4 (
    .d (net160),
    .clk (net1),
    .s (net111),
    .r (net112),
    .q (net161)
  );
  dffsr_cell flop7 (
    .d (net162),
    .clk (net1),
    .s (net111),
    .r (net112),
    .q (net163)
  );
  dffsr_cell flop8 (
    .d (net164),
    .clk (net1),
    .s (net111),
    .r (net112),
    .q (net165)
  );
  dffsr_cell flop9 (
    .d (net166),
    .clk (net1),
    .s (net167),
    .r (net168),
    .q (net44),
    .notq (net169)
  );
  mux_cell mux4 (
    .a (net44),
    .b (net169),
    .sel (net170),
    .out (net171)
  );
  xor_cell xor4 (
    .a (net53),
    .b (net171),
    .out (net172)
  );
  dffsr_cell flop10 (
    .d (net173),
    .clk (net1),
    .s (net168),
    .r (net167),
    .q (net53),
    .notq (net174)
  );
  and_cell and31 (
    .a (net44),
    .b (net53),
    .out (net175)
  );
  and_cell and32 (
    .a (net174),
    .b (net169),
    .out (net176)
  );
  mux_cell mux5 (
    .a (net175),
    .b (net176),
    .sel (net170),
    .out (net177)
  );
  xor_cell xor5 (
    .a (net61),
    .b (net177),
    .out (net178)
  );
  dffsr_cell flop20 (
    .d (net179),
    .clk (net1),
    .s (net168),
    .r (net167),
    .q (net61),
    .notq (net180)
  );
  and_cell and33 (
    .a (net175),
    .b (net61),
    .out (net181)
  );
  and_cell and34 (
    .a (net180),
    .b (net176),
    .out (net182)
  );
  mux_cell mux6 (
    .a (net181),
    .b (net182),
    .sel (net170),
    .out (net183)
  );
  xor_cell xor6 (
    .a (net69),
    .b (net183),
    .out (net184)
  );
  dffsr_cell flop21 (
    .d (net185),
    .clk (net1),
    .s (net167),
    .r (net168),
    .q (net69),
    .notq (net186)
  );
  not_cell not3 (
    .in (net137),
    .out (net167)
  );
  and_cell and35 (
    .a (net187),
    .b (net188),
    .out (net189)
  );
  and_cell and36 (
    .a (net61),
    .b (net69),
    .out (net190)
  );
  and_cell and37 (
    .a (net53),
    .b (net190),
    .out (net191)
  );
  and_cell and38 (
    .a (net192),
    .b (net191),
    .out (net193)
  );
  nand_cell nand1 (
    .a (net44),
    .b (net193),
    .out (net187)
  );
  not_cell not4 (
    .in (net170),
    .out (net192)
  );
  nand_cell nand2 (
    .a (net169),
    .b (net194),
    .out (net188)
  );
  and_cell and39 (
    .a (net170),
    .b (net195),
    .out (net194)
  );
  and_cell and40 (
    .a (net174),
    .b (net196),
    .out (net195)
  );
  and_cell and41 (
    .a (net61),
    .b (net186),
    .out (net196)
  );
  and_cell and42 (
    .a (net189),
    .b (net197),
    .out (net198)
  );
  or_cell or19 (
    .a (net159),
    .b (net161),
    .out (net199)
  );
  nand_cell nand3 (
    .a (net159),
    .b (net161),
    .out (net200)
  );
  and_cell and43 (
    .a (net199),
    .b (net200),
    .out (net201)
  );
  and_cell and44 (
    .a (net201),
    .b (net26),
    .out (net197)
  );
  and_cell and45 (
    .a (net202),
    .b (net161),
    .out (net170)
  );
  not_cell not5 (
    .in (net159),
    .out (net202)
  );
  dffsr_cell flop22 (
    .d (net203),
    .clk (net1),
    .s (net204),
    .r (net205),
    .q (net77),
    .notq (net206)
  );
  mux_cell mux7 (
    .a (net77),
    .b (net206),
    .sel (net207),
    .out (net208)
  );
  xor_cell xor7 (
    .a (net84),
    .b (net208),
    .out (net209)
  );
  dffsr_cell flop23 (
    .d (net210),
    .clk (net1),
    .s (net204),
    .r (net205),
    .q (net84),
    .notq (net211)
  );
  and_cell and46 (
    .a (net77),
    .b (net84),
    .out (net212)
  );
  and_cell and47 (
    .a (net211),
    .b (net206),
    .out (net213)
  );
  mux_cell mux8 (
    .a (net212),
    .b (net213),
    .sel (net207),
    .out (net214)
  );
  xor_cell xor8 (
    .a (net91),
    .b (net214),
    .out (net215)
  );
  dffsr_cell flop24 (
    .d (net216),
    .clk (net1),
    .s (net204),
    .r (net205),
    .q (net91),
    .notq (net217)
  );
  and_cell and48 (
    .a (net212),
    .b (net91),
    .out (net218)
  );
  and_cell and49 (
    .a (net217),
    .b (net213),
    .out (net219)
  );
  mux_cell mux9 (
    .a (net218),
    .b (net219),
    .sel (net207),
    .out (net220)
  );
  xor_cell xor9 (
    .a (net98),
    .b (net220),
    .out (net221)
  );
  dffsr_cell flop25 (
    .d (net222),
    .clk (net1),
    .s (net205),
    .r (net204),
    .q (net98),
    .notq (net223)
  );
  not_cell not6 (
    .in (net137),
    .out (net204)
  );
  and_cell and50 (
    .a (net224),
    .b (net225),
    .out (net226)
  );
  nand_cell nand4 (
    .a (net77),
    .b (net227),
    .out (net224)
  );
  nand_cell nand5 (
    .a (net206),
    .b (net228),
    .out (net225)
  );
  and_cell and59 (
    .a (net226),
    .b (net229),
    .out (net230)
  );
  or_cell or20 (
    .a (net165),
    .b (net163),
    .out (net231)
  );
  nand_cell nand6 (
    .a (net165),
    .b (net163),
    .out (net232)
  );
  and_cell and60 (
    .a (net231),
    .b (net232),
    .out (net233)
  );
  and_cell and61 (
    .a (net233),
    .b (net26),
    .out (net229)
  );
  and_cell and62 (
    .a (net234),
    .b (net163),
    .out (net207)
  );
  not_cell not8 (
    .in (net165),
    .out (net234)
  );
  dffsr_cell flop15 (
    .d (net235),
    .clk (net1),
    .s (net236),
    .r (net237),
    .q (net75),
    .notq (net238)
  );
  mux_cell mux10 (
    .a (net75),
    .b (net238),
    .sel (net239),
    .out (net240)
  );
  xor_cell xor10 (
    .a (net82),
    .b (net240),
    .out (net241)
  );
  dffsr_cell flop16 (
    .d (net242),
    .clk (net1),
    .s (net236),
    .r (net237),
    .q (net82),
    .notq (net243)
  );
  and_cell and51 (
    .a (net75),
    .b (net82),
    .out (net244)
  );
  and_cell and52 (
    .a (net243),
    .b (net238),
    .out (net245)
  );
  mux_cell mux11 (
    .a (net244),
    .b (net245),
    .sel (net239),
    .out (net246)
  );
  xor_cell xor11 (
    .a (net89),
    .b (net246),
    .out (net247)
  );
  dffsr_cell flop17 (
    .d (net248),
    .clk (net1),
    .s (net236),
    .r (net237),
    .q (net89),
    .notq (net249)
  );
  and_cell and53 (
    .a (net244),
    .b (net89),
    .out (net250)
  );
  and_cell and54 (
    .a (net249),
    .b (net245),
    .out (net251)
  );
  mux_cell mux12 (
    .a (net250),
    .b (net251),
    .sel (net239),
    .out (net252)
  );
  xor_cell xor12 (
    .a (net96),
    .b (net252),
    .out (net253)
  );
  dffsr_cell flop28 (
    .d (net254),
    .clk (net1),
    .s (net236),
    .r (net237),
    .q (net96),
    .notq (net255)
  );
  not_cell not7 (
    .in (net137),
    .out (net237)
  );
  and_cell and57 (
    .a (net256),
    .b (net257),
    .out (net258)
  );
  nand_cell nand10 (
    .a (net75),
    .b (net259),
    .out (net256)
  );
  nand_cell nand11 (
    .a (net238),
    .b (net260),
    .out (net257)
  );
  and_cell and58 (
    .a (net258),
    .b (net261),
    .out (net262)
  );
  or_cell or21 (
    .a (net157),
    .b (net155),
    .out (net263)
  );
  nand_cell nand12 (
    .a (net157),
    .b (net155),
    .out (net264)
  );
  and_cell and66 (
    .a (net263),
    .b (net264),
    .out (net265)
  );
  and_cell and82 (
    .a (net265),
    .b (net26),
    .out (net261)
  );
  and_cell and83 (
    .a (net266),
    .b (net155),
    .out (net239)
  );
  not_cell not10 (
    .in (net157),
    .out (net266)
  );
  and_cell and84 (
    .a (net218),
    .b (net98),
    .out (net267)
  );
  and_cell and85 (
    .a (net223),
    .b (net219),
    .out (net268)
  );
  mux_cell mux13 (
    .a (net267),
    .b (net268),
    .sel (net207),
    .out (net269)
  );
  xor_cell xor13 (
    .a (net105),
    .b (net269),
    .out (net270)
  );
  dffsr_cell flop29 (
    .d (net271),
    .clk (net1),
    .s (net204),
    .r (net205),
    .q (net105),
    .notq (net272)
  );
  and_cell and86 (
    .a (net273),
    .b (net274),
    .out (net227)
  );
  and_cell and87 (
    .a (net84),
    .b (net275),
    .out (net274)
  );
  and_cell and88 (
    .a (net91),
    .b (net276),
    .out (net275)
  );
  and_cell and89 (
    .a (net277),
    .b (net105),
    .out (net276)
  );
  not_cell not11 (
    .in (net98),
    .out (net277)
  );
  not_cell not12 (
    .in (net207),
    .out (net273)
  );
  and_cell and90 (
    .a (net207),
    .b (net278),
    .out (net228)
  );
  and_cell and91 (
    .a (net211),
    .b (net279),
    .out (net278)
  );
  and_cell and92 (
    .a (net91),
    .b (net280),
    .out (net279)
  );
  and_cell and93 (
    .a (net98),
    .b (net272),
    .out (net280)
  );
  and_cell and94 (
    .a (net281),
    .b (net282),
    .out (net259)
  );
  not_cell not13 (
    .in (net239),
    .out (net281)
  );
  and_cell and95 (
    .a (net283),
    .b (net239),
    .out (net260)
  );
  and_cell and96 (
    .a (net82),
    .b (net284),
    .out (net282)
  );
  and_cell and97 (
    .a (net249),
    .b (net96),
    .out (net284)
  );
  and_cell and98 (
    .a (net249),
    .b (net255),
    .out (net285)
  );
  and_cell and99 (
    .a (net243),
    .b (net285),
    .out (net283)
  );
  and_cell and100 (
    .a (net41),
    .b (net286),
    .out (net287)
  );
  and_cell and101 (
    .a (net40),
    .b (net286),
    .out (net288)
  );
  and_cell and102 (
    .a (net46),
    .b (net289),
    .out (net290)
  );
  or_cell or22 (
    .a (net287),
    .b (net288),
    .out (net291)
  );
  or_cell or23 (
    .a (net291),
    .b (net290),
    .out (net292)
  );
  dffsr_cell flop33 (
    .d (net293),
    .clk (net1),
    .s (net294),
    .r (net295),
    .q (net47),
    .notq (net296)
  );
  mux_cell mux14 (
    .a (net47),
    .b (net296),
    .sel (net297),
    .out (net298)
  );
  xor_cell xor14 (
    .a (net55),
    .b (net298),
    .out (net299)
  );
  dffsr_cell flop34 (
    .d (net300),
    .clk (net1),
    .s (net294),
    .r (net295),
    .q (net55),
    .notq (net301)
  );
  and_cell and103 (
    .a (net47),
    .b (net55),
    .out (net302)
  );
  and_cell and104 (
    .a (net301),
    .b (net296),
    .out (net303)
  );
  mux_cell mux15 (
    .a (net302),
    .b (net303),
    .sel (net297),
    .out (net304)
  );
  xor_cell xor15 (
    .a (net63),
    .b (net304),
    .out (net305)
  );
  dffsr_cell flop35 (
    .d (net306),
    .clk (net1),
    .s (net294),
    .r (net295),
    .q (net63),
    .notq (net307)
  );
  and_cell and105 (
    .a (net302),
    .b (net63),
    .out (net308)
  );
  and_cell and106 (
    .a (net307),
    .b (net303),
    .out (net309)
  );
  mux_cell mux16 (
    .a (net308),
    .b (net309),
    .sel (net297),
    .out (net310)
  );
  xor_cell xor16 (
    .a (net71),
    .b (net310),
    .out (net311)
  );
  dffsr_cell flop36 (
    .d (net312),
    .clk (net1),
    .s (net294),
    .r (net295),
    .q (net71),
    .notq (net313)
  );
  dffsr_cell flop37 (
    .d (net314),
    .clk (net1),
    .s (net315),
    .r (net316),
    .q (net79),
    .notq (net317)
  );
  mux_cell mux17 (
    .a (net79),
    .b (net317),
    .sel (net318),
    .out (net319)
  );
  xor_cell xor17 (
    .a (net86),
    .b (net319),
    .out (net320)
  );
  dffsr_cell flop38 (
    .d (net321),
    .clk (net1),
    .s (net322),
    .r (net323),
    .q (net86),
    .notq (net324)
  );
  and_cell and107 (
    .a (net79),
    .b (net86),
    .out (net325)
  );
  and_cell and108 (
    .a (net324),
    .b (net317),
    .out (net326)
  );
  mux_cell mux18 (
    .a (net325),
    .b (net326),
    .sel (net318),
    .out (net327)
  );
  xor_cell xor18 (
    .a (net93),
    .b (net327),
    .out (net328)
  );
  dffsr_cell flop39 (
    .d (net329),
    .clk (net1),
    .s (net330),
    .r (net331),
    .q (net93),
    .notq (net332)
  );
  and_cell and109 (
    .a (net325),
    .b (net93),
    .out (net333)
  );
  and_cell and110 (
    .a (net332),
    .b (net326),
    .out (net334)
  );
  mux_cell mux19 (
    .a (net333),
    .b (net334),
    .sel (net318),
    .out (net335)
  );
  xor_cell xor19 (
    .a (net100),
    .b (net335),
    .out (net336)
  );
  dffsr_cell flop40 (
    .d (net337),
    .clk (net1),
    .s (net338),
    .r (net339),
    .q (net100),
    .notq (net340)
  );
  and_cell and111 (
    .a (net333),
    .b (net100),
    .out (net341)
  );
  and_cell and112 (
    .a (net340),
    .b (net334),
    .out (net342)
  );
  mux_cell mux20 (
    .a (net341),
    .b (net342),
    .sel (net318),
    .out (net343)
  );
  xor_cell xor20 (
    .a (net107),
    .b (net343),
    .out (net344)
  );
  dffsr_cell flop41 (
    .d (net345),
    .clk (net1),
    .s (net339),
    .r (net338),
    .q (net107),
    .notq (net346)
  );
  and_cell and113 (
    .a (net63),
    .b (net71),
    .out (net347)
  );
  and_cell and114 (
    .a (net55),
    .b (net347),
    .out (net348)
  );
  and_cell and117 (
    .a (net301),
    .b (net349),
    .out (net350)
  );
  and_cell and118 (
    .a (net307),
    .b (net313),
    .out (net349)
  );
  xor_cell xor22 (
    .a (net351),
    .b (net352),
    .out (net353)
  );
  not_cell not14 (
    .in (net353),
    .out (net354)
  );
  and_cell and116 (
    .a (net47),
    .b (net348),
    .out (net352)
  );
  nand_cell nand13 (
    .a (net296),
    .b (net350),
    .out (net351)
  );
  and_cell and115 (
    .a (net354),
    .b (net355),
    .out (net356)
  );
  or_cell or24 (
    .a (net352),
    .b (net351),
    .out (net357)
  );
  and_cell and119 (
    .a (net357),
    .b (net354),
    .out (net358)
  );
  not_cell not18 (
    .in (net357),
    .out (net355)
  );
  or_cell or25 (
    .a (net356),
    .b (net295),
    .out (net359)
  );
  not_cell not19 (
    .in (net137),
    .out (net295)
  );
  dffsr_cell flop44 (
    .d (net360),
    .clk (net338),
    .s (net361),
    .r (net361),
    .q (net362),
    .notq (net360)
  );
  not_cell not20 (
    .in (net137),
    .out (net338)
  );
  and_cell and120 (
    .a (net362),
    .b (net338),
    .out (net315)
  );
  and_cell and121 (
    .a (net338),
    .b (net360),
    .out (net316)
  );
  and_cell and122 (
    .a (net362),
    .b (net338),
    .out (net322)
  );
  and_cell and123 (
    .a (net338),
    .b (net360),
    .out (net323)
  );
  and_cell and124 (
    .a (net362),
    .b (net338),
    .out (net331)
  );
  and_cell and125 (
    .a (net338),
    .b (net360),
    .out (net330)
  );
  and_cell and126 (
    .a (net79),
    .b (net363),
    .out (net17)
  );
  and_cell and127 (
    .a (net317),
    .b (net364),
    .out (net16)
  );
  and_cell and128 (
    .a (net93),
    .b (net365),
    .out (net366)
  );
  and_cell and129 (
    .a (net332),
    .b (net367),
    .out (net368)
  );
  and_cell and130 (
    .a (net86),
    .b (net366),
    .out (net363)
  );
  and_cell and131 (
    .a (net324),
    .b (net368),
    .out (net364)
  );
  and_cell and132 (
    .a (net340),
    .b (net107),
    .out (net365)
  );
  and_cell and133 (
    .a (net340),
    .b (net346),
    .out (net367)
  );
  and_cell and138 (
    .a (net338),
    .b (net360),
    .out (net369)
  );
  and_cell and139 (
    .a (net362),
    .b (net338),
    .out (net370)
  );
  and_cell and135 (
    .a (net371),
    .b (net2),
    .out (net137)
  );
  or_cell or26 (
    .a (net17),
    .b (net16),
    .out (net372)
  );
  not_cell not22 (
    .in (net373),
    .out (net371)
  );
  not_cell not21 (
    .in (net2),
    .out (net112)
  );
  xor_cell xor25 (
    .a (net100),
    .b (net98),
    .out (net374)
  );
  not_cell not9 (
    .in (net374),
    .out (net375)
  );
  xor_cell xor26 (
    .a (net93),
    .b (net91),
    .out (net376)
  );
  not_cell not23 (
    .in (net376),
    .out (net377)
  );
  xor_cell xor27 (
    .a (net86),
    .b (net84),
    .out (net378)
  );
  not_cell not24 (
    .in (net378),
    .out (net379)
  );
  xor_cell xor28 (
    .a (net79),
    .b (net77),
    .out (net380)
  );
  not_cell not25 (
    .in (net380),
    .out (net381)
  );
  xor_cell xor34 (
    .a (net107),
    .b (net105),
    .out (net382)
  );
  not_cell not31 (
    .in (net382),
    .out (net383)
  );
  and_cell and65 (
    .a (net375),
    .b (net383),
    .out (net384)
  );
  and_cell and134 (
    .a (net379),
    .b (net377),
    .out (net385)
  );
  and_cell and137 (
    .a (net381),
    .b (net385),
    .out (net386)
  );
  and_cell and140 (
    .a (net386),
    .b (net384),
    .out (net387)
  );
  xor_cell xor29 (
    .a (net100),
    .b (net96),
    .out (net388)
  );
  not_cell not26 (
    .in (net388),
    .out (net389)
  );
  xor_cell xor30 (
    .a (net93),
    .b (net89),
    .out (net390)
  );
  not_cell not27 (
    .in (net390),
    .out (net391)
  );
  xor_cell xor31 (
    .a (net86),
    .b (net82),
    .out (net392)
  );
  not_cell not28 (
    .in (net392),
    .out (net393)
  );
  xor_cell xor32 (
    .a (net79),
    .b (net75),
    .out (net394)
  );
  not_cell not29 (
    .in (net394),
    .out (net395)
  );
  xor_cell xor33 (
    .a (net107),
    .b (net396),
    .out (net397)
  );
  not_cell not30 (
    .in (net397),
    .out (net398)
  );
  and_cell and141 (
    .a (net389),
    .b (net398),
    .out (net399)
  );
  and_cell and142 (
    .a (net393),
    .b (net391),
    .out (net400)
  );
  and_cell and143 (
    .a (net395),
    .b (net400),
    .out (net401)
  );
  and_cell and144 (
    .a (net401),
    .b (net399),
    .out (net402)
  );
  or_cell or28 (
    .a (net403),
    .b (net370),
    .out (net404)
  );
  or_cell or29 (
    .a (net369),
    .b (net405),
    .out (net406)
  );
  xor_cell xor36 (
    .a (net47),
    .b (net407),
    .out (net408)
  );
  not_cell not32 (
    .in (net408),
    .out (net409)
  );
  xor_cell xor37 (
    .a (net55),
    .b (net410),
    .out (net411)
  );
  not_cell not33 (
    .in (net411),
    .out (net412)
  );
  and_cell and145 (
    .a (net409),
    .b (net412),
    .out (net413)
  );
  xor_cell xor38 (
    .a (net63),
    .b (net414),
    .out (net415)
  );
  not_cell not34 (
    .in (net415),
    .out (net416)
  );
  xor_cell xor39 (
    .a (net71),
    .b (net417),
    .out (net418)
  );
  not_cell not35 (
    .in (net418),
    .out (net419)
  );
  and_cell and146 (
    .a (net416),
    .b (net419),
    .out (net420)
  );
  and_cell and147 (
    .a (net413),
    .b (net420),
    .out (net421)
  );
  xor_cell xor35 (
    .a (net422),
    .b (net422),
    .out (net423)
  );
  xor_cell xor40 (
    .a (net42),
    .b (net423),
    .out (net424)
  );
  and_cell and149 (
    .a (net423),
    .b (net42),
    .out (net425)
  );
  xor_cell xor41 (
    .a (net422),
    .b (net424),
    .out (net407)
  );
  and_cell and148 (
    .a (net424),
    .b (net422),
    .out (net426)
  );
  or_cell or31 (
    .a (net425),
    .b (net426),
    .out (net427)
  );
  xor_cell xor42 (
    .a (net422),
    .b (net422),
    .out (net428)
  );
  xor_cell xor43 (
    .a (net51),
    .b (net428),
    .out (net429)
  );
  and_cell and150 (
    .a (net428),
    .b (net51),
    .out (net430)
  );
  xor_cell xor44 (
    .a (net427),
    .b (net429),
    .out (net410)
  );
  and_cell and151 (
    .a (net429),
    .b (net427),
    .out (net431)
  );
  or_cell or32 (
    .a (net430),
    .b (net431),
    .out (net432)
  );
  xor_cell xor45 (
    .a (net422),
    .b (net433),
    .out (net434)
  );
  xor_cell xor46 (
    .a (net59),
    .b (net434),
    .out (net435)
  );
  and_cell and152 (
    .a (net434),
    .b (net59),
    .out (net436)
  );
  xor_cell xor47 (
    .a (net432),
    .b (net435),
    .out (net414)
  );
  and_cell and153 (
    .a (net435),
    .b (net432),
    .out (net437)
  );
  or_cell or33 (
    .a (net436),
    .b (net437),
    .out (net438)
  );
  xor_cell xor48 (
    .a (net422),
    .b (net433),
    .out (net439)
  );
  xor_cell xor49 (
    .a (net67),
    .b (net439),
    .out (net440)
  );
  xor_cell xor50 (
    .a (net438),
    .b (net440),
    .out (net417)
  );
  xor_cell xor51 (
    .a (net47),
    .b (net441),
    .out (net442)
  );
  not_cell not36 (
    .in (net442),
    .out (net443)
  );
  xor_cell xor52 (
    .a (net55),
    .b (net444),
    .out (net445)
  );
  not_cell not37 (
    .in (net445),
    .out (net446)
  );
  and_cell and155 (
    .a (net443),
    .b (net446),
    .out (net447)
  );
  xor_cell xor53 (
    .a (net63),
    .b (net448),
    .out (net449)
  );
  not_cell not38 (
    .in (net449),
    .out (net450)
  );
  xor_cell xor54 (
    .a (net71),
    .b (net451),
    .out (net452)
  );
  not_cell not39 (
    .in (net452),
    .out (net453)
  );
  and_cell and156 (
    .a (net450),
    .b (net453),
    .out (net454)
  );
  and_cell and157 (
    .a (net447),
    .b (net454),
    .out (net455)
  );
  xor_cell xor55 (
    .a (net456),
    .b (net457),
    .out (net458)
  );
  xor_cell xor56 (
    .a (net42),
    .b (net458),
    .out (net459)
  );
  and_cell and158 (
    .a (net458),
    .b (net42),
    .out (net460)
  );
  xor_cell xor57 (
    .a (net456),
    .b (net459),
    .out (net441)
  );
  and_cell and159 (
    .a (net459),
    .b (net456),
    .out (net461)
  );
  or_cell or34 (
    .a (net460),
    .b (net461),
    .out (net462)
  );
  xor_cell xor58 (
    .a (net456),
    .b (net456),
    .out (net463)
  );
  xor_cell xor59 (
    .a (net51),
    .b (net463),
    .out (net464)
  );
  and_cell and160 (
    .a (net463),
    .b (net51),
    .out (net465)
  );
  xor_cell xor60 (
    .a (net462),
    .b (net464),
    .out (net444)
  );
  and_cell and161 (
    .a (net464),
    .b (net462),
    .out (net466)
  );
  or_cell or35 (
    .a (net465),
    .b (net466),
    .out (net467)
  );
  xor_cell xor61 (
    .a (net456),
    .b (net457),
    .out (net468)
  );
  xor_cell xor62 (
    .a (net59),
    .b (net468),
    .out (net469)
  );
  and_cell and162 (
    .a (net468),
    .b (net59),
    .out (net470)
  );
  xor_cell xor63 (
    .a (net467),
    .b (net469),
    .out (net448)
  );
  and_cell and163 (
    .a (net469),
    .b (net467),
    .out (net471)
  );
  or_cell or36 (
    .a (net470),
    .b (net471),
    .out (net472)
  );
  xor_cell xor64 (
    .a (net456),
    .b (net457),
    .out (net473)
  );
  xor_cell xor65 (
    .a (net67),
    .b (net473),
    .out (net474)
  );
  xor_cell xor66 (
    .a (net472),
    .b (net474),
    .out (net451)
  );
  xor_cell xor67 (
    .a (net47),
    .b (net475),
    .out (net476)
  );
  not_cell not40 (
    .in (net476),
    .out (net477)
  );
  xor_cell xor68 (
    .a (net55),
    .b (net478),
    .out (net479)
  );
  not_cell not41 (
    .in (net479),
    .out (net480)
  );
  and_cell and154 (
    .a (net477),
    .b (net480),
    .out (net481)
  );
  xor_cell xor69 (
    .a (net63),
    .b (net482),
    .out (net483)
  );
  not_cell not42 (
    .in (net483),
    .out (net484)
  );
  xor_cell xor70 (
    .a (net71),
    .b (net485),
    .out (net486)
  );
  not_cell not43 (
    .in (net486),
    .out (net487)
  );
  and_cell and164 (
    .a (net484),
    .b (net487),
    .out (net488)
  );
  and_cell and165 (
    .a (net481),
    .b (net488),
    .out (net489)
  );
  xor_cell xor71 (
    .a (net490),
    .b (net490),
    .out (net491)
  );
  xor_cell xor72 (
    .a (net42),
    .b (net491),
    .out (net492)
  );
  and_cell and166 (
    .a (net491),
    .b (net42),
    .out (net493)
  );
  xor_cell xor73 (
    .a (net490),
    .b (net492),
    .out (net475)
  );
  and_cell and167 (
    .a (net492),
    .b (net490),
    .out (net494)
  );
  or_cell or37 (
    .a (net493),
    .b (net494),
    .out (net495)
  );
  xor_cell xor74 (
    .a (net490),
    .b (net496),
    .out (net497)
  );
  xor_cell xor75 (
    .a (net51),
    .b (net497),
    .out (net498)
  );
  and_cell and168 (
    .a (net497),
    .b (net51),
    .out (net499)
  );
  xor_cell xor76 (
    .a (net495),
    .b (net498),
    .out (net478)
  );
  and_cell and169 (
    .a (net498),
    .b (net495),
    .out (net500)
  );
  or_cell or38 (
    .a (net499),
    .b (net500),
    .out (net501)
  );
  xor_cell xor77 (
    .a (net490),
    .b (net496),
    .out (net502)
  );
  xor_cell xor78 (
    .a (net59),
    .b (net502),
    .out (net503)
  );
  and_cell and170 (
    .a (net502),
    .b (net59),
    .out (net504)
  );
  xor_cell xor79 (
    .a (net501),
    .b (net503),
    .out (net482)
  );
  and_cell and171 (
    .a (net503),
    .b (net501),
    .out (net505)
  );
  or_cell or39 (
    .a (net504),
    .b (net505),
    .out (net506)
  );
  xor_cell xor80 (
    .a (net490),
    .b (net496),
    .out (net507)
  );
  xor_cell xor81 (
    .a (net67),
    .b (net507),
    .out (net508)
  );
  xor_cell xor82 (
    .a (net506),
    .b (net508),
    .out (net485)
  );
  or_cell or40 (
    .a (net455),
    .b (net509),
    .out (net510)
  );
  xor_cell xor83 (
    .a (net47),
    .b (net511),
    .out (net512)
  );
  not_cell not44 (
    .in (net512),
    .out (net513)
  );
  xor_cell xor84 (
    .a (net55),
    .b (net514),
    .out (net515)
  );
  not_cell not45 (
    .in (net515),
    .out (net516)
  );
  and_cell and172 (
    .a (net513),
    .b (net516),
    .out (net517)
  );
  xor_cell xor85 (
    .a (net63),
    .b (net518),
    .out (net519)
  );
  not_cell not46 (
    .in (net519),
    .out (net520)
  );
  xor_cell xor86 (
    .a (net71),
    .b (net521),
    .out (net522)
  );
  not_cell not47 (
    .in (net522),
    .out (net523)
  );
  and_cell and173 (
    .a (net520),
    .b (net523),
    .out (net524)
  );
  and_cell and174 (
    .a (net517),
    .b (net524),
    .out (net525)
  );
  xor_cell xor87 (
    .a (net526),
    .b (net527),
    .out (net528)
  );
  xor_cell xor88 (
    .a (net44),
    .b (net528),
    .out (net529)
  );
  and_cell and175 (
    .a (net528),
    .b (net44),
    .out (net530)
  );
  xor_cell xor89 (
    .a (net526),
    .b (net529),
    .out (net511)
  );
  and_cell and176 (
    .a (net529),
    .b (net526),
    .out (net531)
  );
  or_cell or41 (
    .a (net530),
    .b (net531),
    .out (net532)
  );
  xor_cell xor90 (
    .a (net526),
    .b (net526),
    .out (net533)
  );
  xor_cell xor91 (
    .a (net53),
    .b (net533),
    .out (net534)
  );
  and_cell and177 (
    .a (net533),
    .b (net53),
    .out (net535)
  );
  xor_cell xor92 (
    .a (net532),
    .b (net534),
    .out (net514)
  );
  and_cell and178 (
    .a (net534),
    .b (net532),
    .out (net536)
  );
  or_cell or42 (
    .a (net535),
    .b (net536),
    .out (net537)
  );
  xor_cell xor93 (
    .a (net526),
    .b (net527),
    .out (net538)
  );
  xor_cell xor94 (
    .a (net61),
    .b (net538),
    .out (net539)
  );
  and_cell and179 (
    .a (net538),
    .b (net61),
    .out (net540)
  );
  xor_cell xor95 (
    .a (net537),
    .b (net539),
    .out (net518)
  );
  and_cell and180 (
    .a (net539),
    .b (net537),
    .out (net541)
  );
  or_cell or43 (
    .a (net540),
    .b (net541),
    .out (net542)
  );
  xor_cell xor96 (
    .a (net526),
    .b (net527),
    .out (net543)
  );
  xor_cell xor97 (
    .a (net69),
    .b (net543),
    .out (net544)
  );
  xor_cell xor98 (
    .a (net542),
    .b (net544),
    .out (net521)
  );
  xor_cell xor99 (
    .a (net47),
    .b (net545),
    .out (net546)
  );
  not_cell not48 (
    .in (net546),
    .out (net547)
  );
  xor_cell xor100 (
    .a (net55),
    .b (net548),
    .out (net549)
  );
  not_cell not49 (
    .in (net549),
    .out (net550)
  );
  and_cell and181 (
    .a (net547),
    .b (net550),
    .out (net551)
  );
  xor_cell xor101 (
    .a (net63),
    .b (net552),
    .out (net553)
  );
  not_cell not50 (
    .in (net553),
    .out (net554)
  );
  xor_cell xor102 (
    .a (net71),
    .b (net555),
    .out (net556)
  );
  not_cell not51 (
    .in (net556),
    .out (net557)
  );
  and_cell and182 (
    .a (net554),
    .b (net557),
    .out (net558)
  );
  and_cell and183 (
    .a (net551),
    .b (net558),
    .out (net559)
  );
  xor_cell xor103 (
    .a (net560),
    .b (net560),
    .out (net561)
  );
  xor_cell xor104 (
    .a (net44),
    .b (net561),
    .out (net562)
  );
  and_cell and184 (
    .a (net561),
    .b (net44),
    .out (net563)
  );
  xor_cell xor105 (
    .a (net560),
    .b (net562),
    .out (net545)
  );
  and_cell and185 (
    .a (net562),
    .b (net560),
    .out (net564)
  );
  or_cell or44 (
    .a (net563),
    .b (net564),
    .out (net565)
  );
  xor_cell xor106 (
    .a (net560),
    .b (net566),
    .out (net567)
  );
  xor_cell xor107 (
    .a (net53),
    .b (net567),
    .out (net568)
  );
  and_cell and186 (
    .a (net567),
    .b (net53),
    .out (net569)
  );
  xor_cell xor108 (
    .a (net565),
    .b (net568),
    .out (net548)
  );
  and_cell and187 (
    .a (net568),
    .b (net565),
    .out (net570)
  );
  or_cell or45 (
    .a (net569),
    .b (net570),
    .out (net571)
  );
  xor_cell xor109 (
    .a (net560),
    .b (net566),
    .out (net572)
  );
  xor_cell xor110 (
    .a (net61),
    .b (net572),
    .out (net573)
  );
  and_cell and188 (
    .a (net572),
    .b (net61),
    .out (net574)
  );
  xor_cell xor111 (
    .a (net571),
    .b (net573),
    .out (net552)
  );
  and_cell and189 (
    .a (net573),
    .b (net571),
    .out (net575)
  );
  or_cell or46 (
    .a (net574),
    .b (net575),
    .out (net576)
  );
  xor_cell xor112 (
    .a (net560),
    .b (net566),
    .out (net577)
  );
  xor_cell xor113 (
    .a (net69),
    .b (net577),
    .out (net578)
  );
  xor_cell xor114 (
    .a (net576),
    .b (net578),
    .out (net555)
  );
  or_cell or47 (
    .a (net525),
    .b (net579),
    .out (net580)
  );
  xor_cell xor115 (
    .a (net47),
    .b (net581),
    .out (net582)
  );
  not_cell not52 (
    .in (net582),
    .out (net583)
  );
  xor_cell xor116 (
    .a (net55),
    .b (net584),
    .out (net585)
  );
  not_cell not53 (
    .in (net585),
    .out (net586)
  );
  and_cell and190 (
    .a (net583),
    .b (net586),
    .out (net587)
  );
  xor_cell xor117 (
    .a (net63),
    .b (net588),
    .out (net589)
  );
  not_cell not54 (
    .in (net589),
    .out (net590)
  );
  xor_cell xor118 (
    .a (net71),
    .b (net591),
    .out (net592)
  );
  not_cell not55 (
    .in (net592),
    .out (net593)
  );
  and_cell and191 (
    .a (net590),
    .b (net593),
    .out (net594)
  );
  and_cell and192 (
    .a (net587),
    .b (net594),
    .out (net595)
  );
  xor_cell xor119 (
    .a (net596),
    .b (net596),
    .out (net597)
  );
  xor_cell xor120 (
    .a (net44),
    .b (net597),
    .out (net598)
  );
  and_cell and193 (
    .a (net597),
    .b (net44),
    .out (net599)
  );
  xor_cell xor121 (
    .a (net596),
    .b (net598),
    .out (net581)
  );
  and_cell and194 (
    .a (net598),
    .b (net596),
    .out (net600)
  );
  or_cell or48 (
    .a (net599),
    .b (net600),
    .out (net601)
  );
  xor_cell xor122 (
    .a (net596),
    .b (net596),
    .out (net602)
  );
  xor_cell xor123 (
    .a (net53),
    .b (net602),
    .out (net603)
  );
  and_cell and195 (
    .a (net602),
    .b (net53),
    .out (net604)
  );
  xor_cell xor124 (
    .a (net601),
    .b (net603),
    .out (net584)
  );
  and_cell and196 (
    .a (net603),
    .b (net601),
    .out (net605)
  );
  or_cell or49 (
    .a (net604),
    .b (net605),
    .out (net606)
  );
  xor_cell xor125 (
    .a (net596),
    .b (net607),
    .out (net608)
  );
  xor_cell xor126 (
    .a (net61),
    .b (net608),
    .out (net609)
  );
  and_cell and197 (
    .a (net608),
    .b (net61),
    .out (net610)
  );
  xor_cell xor127 (
    .a (net606),
    .b (net609),
    .out (net588)
  );
  and_cell and198 (
    .a (net609),
    .b (net606),
    .out (net611)
  );
  or_cell or50 (
    .a (net610),
    .b (net611),
    .out (net612)
  );
  xor_cell xor128 (
    .a (net596),
    .b (net607),
    .out (net613)
  );
  xor_cell xor129 (
    .a (net69),
    .b (net613),
    .out (net614)
  );
  xor_cell xor130 (
    .a (net612),
    .b (net614),
    .out (net591)
  );
  or_cell or51 (
    .a (net595),
    .b (net580),
    .out (net615)
  );
  or_cell or52 (
    .a (net421),
    .b (net510),
    .out (net616)
  );
  xor_cell xor131 (
    .a (net47),
    .b (net42),
    .out (net617)
  );
  not_cell not56 (
    .in (net617),
    .out (net618)
  );
  xor_cell xor132 (
    .a (net55),
    .b (net51),
    .out (net619)
  );
  not_cell not57 (
    .in (net619),
    .out (net620)
  );
  and_cell and199 (
    .a (net618),
    .b (net620),
    .out (net621)
  );
  xor_cell xor133 (
    .a (net63),
    .b (net59),
    .out (net622)
  );
  not_cell not58 (
    .in (net622),
    .out (net623)
  );
  xor_cell xor134 (
    .a (net71),
    .b (net67),
    .out (net624)
  );
  not_cell not59 (
    .in (net624),
    .out (net625)
  );
  and_cell and200 (
    .a (net623),
    .b (net625),
    .out (net626)
  );
  and_cell and201 (
    .a (net621),
    .b (net626),
    .out (net627)
  );
  xor_cell xor135 (
    .a (net47),
    .b (net44),
    .out (net628)
  );
  not_cell not60 (
    .in (net628),
    .out (net629)
  );
  xor_cell xor136 (
    .a (net55),
    .b (net53),
    .out (net630)
  );
  not_cell not61 (
    .in (net630),
    .out (net631)
  );
  and_cell and202 (
    .a (net629),
    .b (net631),
    .out (net632)
  );
  xor_cell xor137 (
    .a (net63),
    .b (net61),
    .out (net633)
  );
  not_cell not62 (
    .in (net633),
    .out (net634)
  );
  xor_cell xor138 (
    .a (net71),
    .b (net69),
    .out (net635)
  );
  not_cell not63 (
    .in (net635),
    .out (net636)
  );
  and_cell and203 (
    .a (net634),
    .b (net636),
    .out (net637)
  );
  and_cell and204 (
    .a (net632),
    .b (net637),
    .out (net638)
  );
  or_cell or53 (
    .a (net559),
    .b (net638),
    .out (net579)
  );
  or_cell or54 (
    .a (net489),
    .b (net627),
    .out (net509)
  );
  or_cell or55 (
    .a (net402),
    .b (net616),
    .out (net405)
  );
  or_cell or56 (
    .a (net387),
    .b (net615),
    .out (net403)
  );
  dffsr_cell flop30 (
    .d (net372),
    .clk (net1),
    .s (net639),
    .r (net112),
    .q (net373)
  );
  and_cell and205 (
    .a (net66),
    .b (net58),
    .out (net640)
  );
  and_cell and206 (
    .a (net640),
    .b (net50),
    .out (net641)
  );
  and_cell and207 (
    .a (net66),
    .b (net58),
    .out (net642)
  );
  and_cell and208 (
    .a (net642),
    .b (net643),
    .out (net644)
  );
  and_cell and209 (
    .a (net66),
    .b (net645),
    .out (net646)
  );
  and_cell and210 (
    .a (net646),
    .b (net50),
    .out (net647)
  );
  and_cell and211 (
    .a (net66),
    .b (net645),
    .out (net648)
  );
  and_cell and212 (
    .a (net648),
    .b (net643),
    .out (net649)
  );
  and_cell and213 (
    .a (net650),
    .b (net58),
    .out (net651)
  );
  and_cell and214 (
    .a (net651),
    .b (net50),
    .out (net652)
  );
  and_cell and215 (
    .a (net650),
    .b (net58),
    .out (net653)
  );
  and_cell and216 (
    .a (net653),
    .b (net643),
    .out (net654)
  );
  and_cell and217 (
    .a (net650),
    .b (net645),
    .out (net655)
  );
  and_cell and218 (
    .a (net655),
    .b (net50),
    .out (net656)
  );
  and_cell and219 (
    .a (net650),
    .b (net645),
    .out (net657)
  );
  and_cell and220 (
    .a (net657),
    .b (net643),
    .out (net658)
  );
  not_cell not64 (
    .in (net50),
    .out (net643)
  );
  not_cell not65 (
    .in (net58),
    .out (net645)
  );
  not_cell not66 (
    .in (net66),
    .out (net650)
  );
  and_cell and221 (
    .a (net74),
    .b (net641),
    .out (net659)
  );
  and_cell and222 (
    .a (net74),
    .b (net644),
    .out (net660)
  );
  and_cell and223 (
    .a (net74),
    .b (net647),
    .out (net661)
  );
  and_cell and224 (
    .a (net74),
    .b (net649),
    .out (net662)
  );
  and_cell and225 (
    .a (net74),
    .b (net652),
    .out (net663)
  );
  and_cell and226 (
    .a (net74),
    .b (net654),
    .out (net664)
  );
  and_cell and227 (
    .a (net74),
    .b (net656),
    .out (net665)
  );
  and_cell and228 (
    .a (net74),
    .b (net658),
    .out (net666)
  );
  and_cell and229 (
    .a (net66),
    .b (net58),
    .out (net667)
  );
  and_cell and230 (
    .a (net667),
    .b (net50),
    .out (net668)
  );
  and_cell and231 (
    .a (net66),
    .b (net58),
    .out (net669)
  );
  and_cell and232 (
    .a (net669),
    .b (net670),
    .out (net671)
  );
  and_cell and233 (
    .a (net66),
    .b (net672),
    .out (net673)
  );
  and_cell and234 (
    .a (net673),
    .b (net50),
    .out (net674)
  );
  and_cell and235 (
    .a (net66),
    .b (net672),
    .out (net675)
  );
  and_cell and236 (
    .a (net675),
    .b (net670),
    .out (net676)
  );
  and_cell and237 (
    .a (net677),
    .b (net58),
    .out (net678)
  );
  and_cell and238 (
    .a (net678),
    .b (net50),
    .out (net679)
  );
  and_cell and239 (
    .a (net677),
    .b (net58),
    .out (net680)
  );
  and_cell and240 (
    .a (net680),
    .b (net670),
    .out (net681)
  );
  and_cell and241 (
    .a (net677),
    .b (net672),
    .out (net682)
  );
  and_cell and242 (
    .a (net682),
    .b (net50),
    .out (net683)
  );
  and_cell and243 (
    .a (net677),
    .b (net672),
    .out (net684)
  );
  and_cell and244 (
    .a (net684),
    .b (net670),
    .out (net685)
  );
  not_cell not67 (
    .in (net50),
    .out (net670)
  );
  not_cell not68 (
    .in (net58),
    .out (net672)
  );
  not_cell not69 (
    .in (net66),
    .out (net677)
  );
  and_cell and245 (
    .a (net686),
    .b (net668),
    .out (net687)
  );
  and_cell and246 (
    .a (net686),
    .b (net671),
    .out (net688)
  );
  and_cell and247 (
    .a (net686),
    .b (net674),
    .out (net689)
  );
  and_cell and248 (
    .a (net686),
    .b (net676),
    .out (net690)
  );
  and_cell and249 (
    .a (net686),
    .b (net679),
    .out (net691)
  );
  and_cell and250 (
    .a (net686),
    .b (net681),
    .out (net692)
  );
  and_cell and251 (
    .a (net686),
    .b (net683),
    .out (net693)
  );
  and_cell and252 (
    .a (net686),
    .b (net685),
    .out (net694)
  );
  not_cell not76 (
    .in (net74),
    .out (net686)
  );
  and_cell and301 (
    .a (net292),
    .b (net659),
    .out (net695)
  );
  and_cell and302 (
    .a (net292),
    .b (net660),
    .out (net696)
  );
  and_cell and303 (
    .a (net292),
    .b (net661),
    .out (net697)
  );
  and_cell and304 (
    .a (net292),
    .b (net662),
    .out (net698)
  );
  and_cell and305 (
    .a (net292),
    .b (net663),
    .out (net699)
  );
  and_cell and306 (
    .a (net292),
    .b (net664),
    .out (net700)
  );
  and_cell and307 (
    .a (net292),
    .b (net665),
    .out (net701)
  );
  and_cell and308 (
    .a (net292),
    .b (net666),
    .out (net702)
  );
  and_cell and309 (
    .a (net292),
    .b (net687),
    .out (net703)
  );
  and_cell and310 (
    .a (net292),
    .b (net688),
    .out (net704)
  );
  and_cell and311 (
    .a (net292),
    .b (net689),
    .out (net705)
  );
  and_cell and312 (
    .a (net292),
    .b (net690),
    .out (net706)
  );
  and_cell and313 (
    .a (net292),
    .b (net691),
    .out (net707)
  );
  or_cell or60 (
    .a (net660),
    .b (net695),
    .out (net708)
  );
  or_cell or63 (
    .a (net661),
    .b (net695),
    .out (net709)
  );
  or_cell or64 (
    .a (net709),
    .b (net696),
    .out (net710)
  );
  or_cell or66 (
    .a (net662),
    .b (net695),
    .out (net711)
  );
  or_cell or67 (
    .a (net711),
    .b (net696),
    .out (net712)
  );
  or_cell or68 (
    .a (net712),
    .b (net697),
    .out (net713)
  );
  or_cell or69 (
    .a (net663),
    .b (net698),
    .out (net714)
  );
  or_cell or70 (
    .a (net714),
    .b (net696),
    .out (net715)
  );
  or_cell or71 (
    .a (net715),
    .b (net697),
    .out (net716)
  );
  or_cell or72 (
    .a (net664),
    .b (net698),
    .out (net717)
  );
  or_cell or73 (
    .a (net717),
    .b (net699),
    .out (net718)
  );
  or_cell or74 (
    .a (net718),
    .b (net697),
    .out (net719)
  );
  or_cell or75 (
    .a (net665),
    .b (net698),
    .out (net720)
  );
  or_cell or76 (
    .a (net720),
    .b (net699),
    .out (net721)
  );
  or_cell or77 (
    .a (net721),
    .b (net700),
    .out (net722)
  );
  or_cell or78 (
    .a (net666),
    .b (net701),
    .out (net723)
  );
  or_cell or79 (
    .a (net723),
    .b (net699),
    .out (net724)
  );
  or_cell or80 (
    .a (net724),
    .b (net700),
    .out (net725)
  );
  or_cell or81 (
    .a (net687),
    .b (net701),
    .out (net726)
  );
  or_cell or82 (
    .a (net726),
    .b (net702),
    .out (net727)
  );
  or_cell or83 (
    .a (net727),
    .b (net700),
    .out (net728)
  );
  or_cell or84 (
    .a (net688),
    .b (net701),
    .out (net729)
  );
  or_cell or85 (
    .a (net729),
    .b (net702),
    .out (net730)
  );
  or_cell or86 (
    .a (net730),
    .b (net703),
    .out (net731)
  );
  or_cell or87 (
    .a (net689),
    .b (net704),
    .out (net732)
  );
  or_cell or88 (
    .a (net732),
    .b (net702),
    .out (net733)
  );
  or_cell or89 (
    .a (net733),
    .b (net703),
    .out (net734)
  );
  or_cell or90 (
    .a (net690),
    .b (net704),
    .out (net735)
  );
  or_cell or91 (
    .a (net735),
    .b (net705),
    .out (net736)
  );
  or_cell or92 (
    .a (net736),
    .b (net703),
    .out (net737)
  );
  or_cell or93 (
    .a (net691),
    .b (net704),
    .out (net738)
  );
  or_cell or94 (
    .a (net738),
    .b (net705),
    .out (net739)
  );
  or_cell or95 (
    .a (net739),
    .b (net706),
    .out (net740)
  );
  or_cell or96 (
    .a (net692),
    .b (net707),
    .out (net741)
  );
  or_cell or97 (
    .a (net741),
    .b (net705),
    .out (net742)
  );
  or_cell or98 (
    .a (net742),
    .b (net706),
    .out (net743)
  );
  or_cell or99 (
    .a (net693),
    .b (net707),
    .out (net744)
  );
  or_cell or100 (
    .a (net744),
    .b (net706),
    .out (net745)
  );
  or_cell or102 (
    .a (net694),
    .b (net707),
    .out (net746)
  );
  and_cell and253 (
    .a (net641),
    .b (net747),
    .out (net748)
  );
  and_cell and254 (
    .a (net19),
    .b (net749),
    .out (net750)
  );
  or_cell or57 (
    .a (net748),
    .b (net750),
    .out (net751)
  );
  dff_cell flop31 (
    .d (net751),
    .clk (net21),
    .q (net18)
  );
  and_cell and255 (
    .a (net708),
    .b (net747),
    .out (net752)
  );
  and_cell and256 (
    .a (net19),
    .b (net753),
    .out (net754)
  );
  or_cell or58 (
    .a (net752),
    .b (net754),
    .out (net755)
  );
  dff_cell flop48 (
    .d (net755),
    .clk (net21),
    .q (net749)
  );
  and_cell and257 (
    .a (net710),
    .b (net747),
    .out (net756)
  );
  and_cell and258 (
    .a (net19),
    .b (net757),
    .out (net758)
  );
  or_cell or59 (
    .a (net756),
    .b (net758),
    .out (net759)
  );
  dff_cell flop49 (
    .d (net759),
    .clk (net21),
    .q (net753)
  );
  and_cell and259 (
    .a (net713),
    .b (net747),
    .out (net760)
  );
  and_cell and260 (
    .a (net19),
    .b (net761),
    .out (net762)
  );
  or_cell or61 (
    .a (net760),
    .b (net762),
    .out (net763)
  );
  dff_cell flop50 (
    .d (net763),
    .clk (net21),
    .q (net757)
  );
  and_cell and261 (
    .a (net716),
    .b (net747),
    .out (net764)
  );
  and_cell and262 (
    .a (net19),
    .b (net765),
    .out (net766)
  );
  or_cell or62 (
    .a (net764),
    .b (net766),
    .out (net767)
  );
  dff_cell flop51 (
    .d (net767),
    .clk (net21),
    .q (net761)
  );
  and_cell and263 (
    .a (net719),
    .b (net747),
    .out (net768)
  );
  and_cell and264 (
    .a (net19),
    .b (net769),
    .out (net770)
  );
  or_cell or65 (
    .a (net768),
    .b (net770),
    .out (net771)
  );
  dff_cell flop52 (
    .d (net771),
    .clk (net21),
    .q (net765)
  );
  and_cell and265 (
    .a (net722),
    .b (net747),
    .out (net772)
  );
  and_cell and266 (
    .a (net19),
    .b (net773),
    .out (net774)
  );
  or_cell or101 (
    .a (net772),
    .b (net774),
    .out (net775)
  );
  dff_cell flop53 (
    .d (net775),
    .clk (net21),
    .q (net769)
  );
  and_cell and267 (
    .a (net725),
    .b (net747),
    .out (net776)
  );
  and_cell and268 (
    .a (net19),
    .b (net777),
    .out (net778)
  );
  or_cell or103 (
    .a (net776),
    .b (net778),
    .out (net779)
  );
  dff_cell flop54 (
    .d (net779),
    .clk (net21),
    .q (net773)
  );
  and_cell and269 (
    .a (net728),
    .b (net747),
    .out (net780)
  );
  and_cell and270 (
    .a (net19),
    .b (net781),
    .out (net782)
  );
  or_cell or104 (
    .a (net780),
    .b (net782),
    .out (net783)
  );
  dff_cell flop55 (
    .d (net783),
    .clk (net21),
    .q (net777)
  );
  and_cell and271 (
    .a (net731),
    .b (net747),
    .out (net784)
  );
  and_cell and272 (
    .a (net19),
    .b (net785),
    .out (net786)
  );
  or_cell or105 (
    .a (net784),
    .b (net786),
    .out (net787)
  );
  dff_cell flop56 (
    .d (net787),
    .clk (net21),
    .q (net781)
  );
  and_cell and273 (
    .a (net734),
    .b (net747),
    .out (net788)
  );
  and_cell and274 (
    .a (net19),
    .b (net789),
    .out (net790)
  );
  or_cell or106 (
    .a (net788),
    .b (net790),
    .out (net791)
  );
  dff_cell flop57 (
    .d (net791),
    .clk (net21),
    .q (net785)
  );
  and_cell and275 (
    .a (net737),
    .b (net747),
    .out (net792)
  );
  and_cell and276 (
    .a (net19),
    .b (net793),
    .out (net794)
  );
  or_cell or107 (
    .a (net792),
    .b (net794),
    .out (net795)
  );
  dff_cell flop58 (
    .d (net795),
    .clk (net21),
    .q (net789)
  );
  and_cell and277 (
    .a (net740),
    .b (net747),
    .out (net796)
  );
  and_cell and278 (
    .a (net19),
    .b (net797),
    .out (net798)
  );
  or_cell or108 (
    .a (net796),
    .b (net798),
    .out (net799)
  );
  dff_cell flop59 (
    .d (net799),
    .clk (net21),
    .q (net793)
  );
  and_cell and279 (
    .a (net743),
    .b (net747),
    .out (net800)
  );
  and_cell and280 (
    .a (net19),
    .b (net801),
    .out (net802)
  );
  or_cell or109 (
    .a (net800),
    .b (net802),
    .out (net803)
  );
  dff_cell flop60 (
    .d (net803),
    .clk (net21),
    .q (net797)
  );
  and_cell and281 (
    .a (net745),
    .b (net747),
    .out (net804)
  );
  and_cell and282 (
    .a (net19),
    .b (net805),
    .out (net806)
  );
  or_cell or110 (
    .a (net804),
    .b (net806),
    .out (net807)
  );
  dff_cell flop61 (
    .d (net807),
    .clk (net21),
    .q (net801)
  );
  dff_cell flop62 (
    .d (net746),
    .clk (net21),
    .q (net805)
  );
  not_cell not70 (
    .in (net19),
    .out (net747)
  );
  nand_cell nand14 (
    .a (net318),
    .b (net808),
    .out (net809)
  );
  nand_cell nand15 (
    .a (net810),
    .b (net809),
    .out (net318)
  );
  not_cell not71 (
    .in (net404),
    .out (net810)
  );
  not_cell not72 (
    .in (net406),
    .out (net808)
  );
  nand_cell nand16 (
    .a (net297),
    .b (net811),
    .out (net812)
  );
  nand_cell nand17 (
    .a (net813),
    .b (net812),
    .out (net297)
  );
  not_cell not73 (
    .in (net358),
    .out (net813)
  );
  not_cell not74 (
    .in (net359),
    .out (net811)
  );
  mux_cell mux21 (
    .a (net165),
    .b (net10),
    .sel (net30),
    .out (net164)
  );
  mux_cell mux22 (
    .a (net163),
    .b (net9),
    .sel (net30),
    .out (net162)
  );
  mux_cell mux23 (
    .a (net161),
    .b (net8),
    .sel (net30),
    .out (net160)
  );
  mux_cell mux24 (
    .a (net159),
    .b (net7),
    .sel (net30),
    .out (net158)
  );
  mux_cell mux25 (
    .a (net157),
    .b (net6),
    .sel (net30),
    .out (net156)
  );
  mux_cell mux26 (
    .a (net155),
    .b (net5),
    .sel (net30),
    .out (net154)
  );
  mux_cell mux27 (
    .a (net115),
    .b (net4),
    .sel (net30),
    .out (net114)
  );
  mux_cell mux28 (
    .a (net113),
    .b (net3),
    .sel (net30),
    .out (net110)
  );
  mux_cell mux29 (
    .a (net42),
    .b (net119),
    .sel (net149),
    .out (net116)
  );
  mux_cell mux30 (
    .a (net51),
    .b (net122),
    .sel (net149),
    .out (net123)
  );
  mux_cell mux31 (
    .a (net59),
    .b (net128),
    .sel (net149),
    .out (net129)
  );
  mux_cell mux32 (
    .a (net67),
    .b (net134),
    .sel (net149),
    .out (net135)
  );
  mux_cell mux33 (
    .a (net44),
    .b (net169),
    .sel (net198),
    .out (net166)
  );
  mux_cell mux34 (
    .a (net53),
    .b (net172),
    .sel (net198),
    .out (net173)
  );
  mux_cell mux35 (
    .a (net61),
    .b (net178),
    .sel (net198),
    .out (net179)
  );
  mux_cell mux36 (
    .a (net69),
    .b (net184),
    .sel (net198),
    .out (net185)
  );
  mux_cell mux37 (
    .a (net77),
    .b (net206),
    .sel (net230),
    .out (net203)
  );
  mux_cell mux38 (
    .a (net84),
    .b (net209),
    .sel (net230),
    .out (net210)
  );
  mux_cell mux39 (
    .a (net91),
    .b (net215),
    .sel (net230),
    .out (net216)
  );
  mux_cell mux40 (
    .a (net98),
    .b (net221),
    .sel (net230),
    .out (net222)
  );
  mux_cell mux41 (
    .a (net105),
    .b (net270),
    .sel (net230),
    .out (net271)
  );
  mux_cell mux42 (
    .a (net75),
    .b (net238),
    .sel (net262),
    .out (net235)
  );
  mux_cell mux43 (
    .a (net82),
    .b (net241),
    .sel (net262),
    .out (net242)
  );
  mux_cell mux44 (
    .a (net89),
    .b (net247),
    .sel (net262),
    .out (net248)
  );
  mux_cell mux45 (
    .a (net96),
    .b (net253),
    .sel (net262),
    .out (net254)
  );
  mux_cell mux46 (
    .a (net47),
    .b (net296),
    .sel (net28),
    .out (net293)
  );
  mux_cell mux47 (
    .a (net55),
    .b (net299),
    .sel (net28),
    .out (net300)
  );
  mux_cell mux48 (
    .a (net63),
    .b (net305),
    .sel (net28),
    .out (net306)
  );
  mux_cell mux49 (
    .a (net71),
    .b (net311),
    .sel (net28),
    .out (net312)
  );
  mux_cell mux50 (
    .a (net79),
    .b (net317),
    .sel (net28),
    .out (net314)
  );
  mux_cell mux51 (
    .a (net86),
    .b (net320),
    .sel (net28),
    .out (net321)
  );
  mux_cell mux52 (
    .a (net93),
    .b (net328),
    .sel (net28),
    .out (net329)
  );
  mux_cell mux53 (
    .a (net100),
    .b (net336),
    .sel (net28),
    .out (net337)
  );
  mux_cell mux54 (
    .a (net107),
    .b (net344),
    .sel (net28),
    .out (net345)
  );
endmodule
